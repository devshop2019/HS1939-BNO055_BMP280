PK
     �J�Z���sQ  sQ     cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_0":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_1":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_2":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_3":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_4":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_5":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_6":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_7":[],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9":["pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4"],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11":["pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5"],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12":["pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13"],"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13":["pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12"],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_0":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_1":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_2":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_3":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9"],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11"],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_6":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_7":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_8":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_9":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_10":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_11":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13"],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12"],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_14":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_15":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_16":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_17":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_18":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_19":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_20":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_21":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_22":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_23":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_24":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_25":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_26":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_27":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_28":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_29":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_30":[],"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_31":[]},"pin_to_color":{"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_0":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_1":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_2":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_3":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_4":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_5":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_6":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_7":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9":"#ff0000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11":"#000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12":"#0000c8","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13":"#00c800","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_0":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_1":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_2":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_3":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4":"#ff0000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_6":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_7":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_8":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_9":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_10":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_11":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12":"#00c800","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13":"#0000c8","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_14":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_15":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_16":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_17":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_18":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_19":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_20":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_21":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_22":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_23":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_24":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_25":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_26":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_27":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_28":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_29":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_30":"#000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_31":"#000000"},"pin_to_state":{"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_0":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_1":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_2":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_3":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_4":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_5":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_6":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_7":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12":"neutral","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_0":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_1":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_2":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_3":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_6":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_7":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_8":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_9":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_10":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_11":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_14":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_15":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_16":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_17":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_18":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_19":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_20":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_21":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_22":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_23":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_24":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_25":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_26":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_27":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_28":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_29":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_30":"neutral","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_31":"neutral"},"next_color_idx":4,"wires_placed_in_order":[["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4"],["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5"],["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13"],["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12"]],"wires_removed_and_placed_in_order":[[[],[["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4"]]],[[],[["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5"]]],[[],[["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13"]]],[[],[["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_0":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_1":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_2":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_3":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_4":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_5":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_6":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_7":"_","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9":"0000000000000000","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11":"0000000000000001","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12":"0000000000000002","pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13":"0000000000000003","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_0":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_1":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_2":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_3":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4":"0000000000000000","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5":"0000000000000001","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_6":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_7":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_8":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_9":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_10":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_11":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12":"0000000000000003","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13":"0000000000000002","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_14":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_15":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_16":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_17":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_18":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_19":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_20":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_21":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_22":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_23":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_24":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_25":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_26":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_27":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_28":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_29":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_30":"_","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_31":"_"},"component_id_to_pins":{"55b2e155-ea99-4963-899f-87089953b4ad":["0","1","2","3","4","5","6","7","9","11","12","13"],"9e7ee43c-5d99-4739-8c51-7e63844aa012":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4"],"0000000000000001":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5"],"0000000000000002":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13"],"0000000000000003":["pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13","pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000002":"Net 2","0000000000000003":"Net 3"},"all_breadboard_info_list":["6725a34c-4ffa-4ca0-a2e3-40a2e834a759_63_2_True_670_-380_up"],"breadboard_info_list":[],"componentsData":[{"compProperties":{},"position":[686.1642294999999,-192.67681750000008],"typeId":"eea59fab-7716-4d23-b5bc-312fc0fc1b61","componentVersion":1,"instanceId":"55b2e155-ea99-4963-899f-87089953b4ad","orientation":"up","circleData":[[647.5,-130.00000000000003],[662.5,-130.00000000000003],[677.5,-130.00000000000003],[692.5,-130.00000000000003],[707.5,-130.00000000000003],[722.5,-130.00000000000003],[737.5000000000003,-130.00000000000003],[752.5000000000003,-130.00000000000003],[772.5196855000002,-208.30708600000006],[772.5196855000002,-197.20472350000003],[772.5196855000002,-186.57480250000003],[772.5196855000002,-175.9448815]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"version":2,"id":"mpn","label":"mpn","description":"","units":"","type":"string","value":"A000066","displayFormat":"input","showOnComp":false,"isVisibleToUser":false},"manufacturer":{"version":2,"id":"manufacturer","label":"manufacturer","description":"","units":"","type":"string","value":"Arduino","displayFormat":"input","showOnComp":false,"isVisibleToUser":false}},"position":[1146.25,-212.4999999999999],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"9e7ee43c-5d99-4739-8c51-7e63844aa012","orientation":"up","circleData":[[1127.5,-69.99999999999997],[1142.5,-69.99999999999997],[1157.5,-69.99999999999997],[1172.5,-69.99999999999997],[1187.5,-69.99999999999997],[1202.5,-69.99999999999997],[1217.5,-69.99999999999997],[1232.5,-69.99999999999997],[1262.5,-69.99999999999997],[1277.5,-69.99999999999997],[1292.5,-69.99999999999997],[1307.5,-69.99999999999997],[1322.5,-69.99999999999997],[1337.5,-69.99999999999997],[1073.5,-354.9999999999999],[1088.5,-354.9999999999999],[1103.5,-354.9999999999999],[1118.5,-354.9999999999999],[1133.5,-354.9999999999999],[1148.5,-354.9999999999999],[1163.5,-354.9999999999999],[1178.5,-354.9999999999999],[1193.5,-354.9999999999999],[1208.5,-354.9999999999999],[1232.5,-354.9999999999999],[1247.5,-354.9999999999999],[1262.5,-354.9999999999999],[1277.5,-354.9999999999999],[1292.5,-354.9999999999999],[1307.5,-354.9999999999999],[1322.5,-354.9999999999999],[1337.5,-354.9999999999999]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"49ec30fc-3e83-4f7c-8694-f4ff0a9e8844\",\"explorerHtmlId\":\"18544677-dba6-4131-8f8e-1adab501b244\",\"nameHtmlId\":\"b5935bff-0d6c-4207-8aca-6b44fa86b7a9\",\"nameInputHtmlId\":\"653200c5-92e2-41f5-aa4a-dcd308d8ac6a\",\"explorerChildHtmlId\":\"b2370268-acec-4e18-86dd-6c83f5bc8cda\",\"explorerCarrotOpenHtmlId\":\"f5e85388-1748-42e5-8294-4b813e91d5fe\",\"explorerCarrotClosedHtmlId\":\"8ad8f949-83a5-4f0f-b698-73ef7915fcff\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"fc7e945d-bc6a-43e8-961b-a9206f82cf1f\",\"explorerHtmlId\":\"e3911c42-5acc-49bb-b26b-0a15426c0b7f\",\"nameHtmlId\":\"d91e670a-9f21-476a-ab23-18de8a7cccf6\",\"nameInputHtmlId\":\"2b7a8c94-ae4e-4d79-9a29-ddde59eee067\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"934da532-3327-461c-bd7b-07171eea47a6\",\"explorerHtmlId\":\"6a210f3f-f26a-49a5-8f02-a2af4f552acf\",\"nameHtmlId\":\"fd985939-700b-44bc-8e71-ab0d33011eeb\",\"nameInputHtmlId\":\"8898983c-28e5-439c-8d2a-2cfcae417483\",\"code\":\"\"},0,","codeLabelPosition":[1146.25,-369.9999999999999],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-380.00000","left":"591.36090","width":"786.13910","height":"335.00000","x":"591.36090","y":"-380.00000"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#ff0000\",\"startPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9\",\"endPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4\",\"rawStartPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_9\",\"rawEndPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"772.5196855000_-208.3070860000\\\",\\\"925.0000000000_-208.3070860000\\\",\\\"925.0000000000_-40.0000000000\\\",\\\"1187.5000000000_-40.0000000000\\\",\\\"1187.5000000000_-70.0000000000\\\"]}\"}","{\"color\":\"#000000\",\"startPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11\",\"endPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5\",\"rawStartPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_11\",\"rawEndPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_5\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"772.5196855000_-197.2047235000\\\",\\\"902.5000000000_-197.2047235000\\\",\\\"902.5000000000_-25.0000000000\\\",\\\"1202.5000000000_-25.0000000000\\\",\\\"1202.5000000000_-70.0000000000\\\"]}\"}","{\"color\":\"#0000c8\",\"startPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12\",\"endPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13\",\"rawStartPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_12\",\"rawEndPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_13\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"772.5196855000_-186.5748025000\\\",\\\"887.5000000000_-186.5748025000\\\",\\\"887.5000000000_27.5000000000\\\",\\\"1337.5000000000_27.5000000000\\\",\\\"1337.5000000000_-70.0000000000\\\"]}\"}","{\"color\":\"#00c800\",\"startPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13\",\"endPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12\",\"rawStartPinId\":\"pin-type-component_55b2e155-ea99-4963-899f-87089953b4ad_13\",\"rawEndPinId\":\"pin-type-component_9e7ee43c-5d99-4739-8c51-7e63844aa012_12\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"772.5196855000_-175.9448815000\\\",\\\"872.5000000000_-175.9448815000\\\",\\\"872.5000000000_5.0000000000\\\",\\\"1322.5000000000_5.0000000000\\\",\\\"1322.5000000000_-70.0000000000\\\"]}\"}"],"projectDescription":""}PK
     �J�Z               jsons/PK
     �J�Z�haZ       jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"DFRobot BNO055 + BMP280","category":["User Defined"],"id":"eea59fab-7716-4d23-b5bc-312fc0fc1b61","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"707f98a2-ba92-4472-bb4e-3eede8d3998f.png","iconPic":"e96e51a4-2e0a-4cc5-ba63-cf190e1d4d54.png","hasComponentImageSvg":false,"componentImageSvgUrl":"","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"11.30711","numDisplayRows":"9.54038","pins":[{"uniquePinIdString":"0","positionMil":"307.59397,59.17355","isAnchorPin":true,"label":""},{"uniquePinIdString":"1","positionMil":"407.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"2","positionMil":"507.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"3","positionMil":"607.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"4","positionMil":"707.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"5","positionMil":"807.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"6","positionMil":"907.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"7","positionMil":"1007.59397,59.17355","isAnchorPin":false,"label":""},{"uniquePinIdString":"9","positionMil":"1141.05854,581.22079","isAnchorPin":false,"label":""},{"uniquePinIdString":"11","positionMil":"1141.05854,507.20504","isAnchorPin":false,"label":""},{"uniquePinIdString":"12","positionMil":"1141.05854,436.33890","isAnchorPin":false,"label":""},{"uniquePinIdString":"13","positionMil":"1141.05854,365.47276","isAnchorPin":false,"label":""}],"pinType":"wired"},"properties":[],"propertiesV2":[]},{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache","hasComponentImageSvg":false,"componentImageSvgUrl":""}]}PK
     �J�Z               images/PK
     �J�Z[�\� \� /   images/707f98a2-ba92-4472-bb4e-3eede8d3998f.png�PNG

   IHDR  �  X   K��)   	pHYs  �  ��+  ��IDATx����y.��Ms�� r�$H�H�)Q�HI$M����d[^S�d�]{��W>G^��9�����q�%+�
�heYb0I� )�����`0����ܴ]�]��u�����3��nwu�N�_}��_����D�,�l�?N���x�/�+
�o`` o��6^~�e�ٳ����Ǒ�fa`````````�#����W\q6l؀n��y�{�b�
�R)$	�@�2b�D���㪸2��011���Q�={�<��z�)�ܹ���0000000000C�Xą��+�����C<ǚ5kp�m���(�lق��&��iJ�E��X�Ⱈ.Q	ש�b�KHsWW^}�U���?�/�@�g���X5+�G5Q���><���X���Pe��� �k����1σb��\#L}fQ����÷��-�رӉп/~��{��}W]u��۩Z�3If��$<��f����qr�N�>��_��ױo�>�&�SM�-$1$b�}#쿘E�����X(]{��˗�/��"���S���~���'���>��|�3���1��2�� r`�N���*�v"�Ν�����|O?�t�i���#SG]:�Z���ejb��I��.����3	��s��h�N�i���M���12�G�p�#��H��<�Egt,���&
�XT��������g�}=�>�O�I�uuuJ�8�SZf��<��y�޽x�G��o���HsCmm61n�O���]:/���,jMc�����Ǝ�D"n�\�q!�Q�k��m�<8����qt���L�Nue��;���	��D�oxC�yC�����n��?�~��_���p�wb�����(�x�r	Y�W����K/�D�L�/�q���[R��-��-5X��W,�ê�uvX�51JzKD�'	�ˇ��������ă�u7(�&�5!���Ӽ틌���M��8rnG:Fp�s=c8g�����������`� ��o�A�&�S��7n��y��eƏ:��ˀL$�5��_�G��� g:H��mҼjA-V����jeV/�E&���>���2���p0�\�KZ*���p�����\d�M��-���������SC8pz���c6���|:(3�C�W��UJ��}뭷R�wa�1o��E`���'O���~�aj�<�Qg�Ջj�~i��	�5��vq=R	�@�_Q�Y��6��b���u���w( Y�A�_�{���_o�6�n���:}���>6�}6�&���ib_m````````P9��8������?�cj�Q__���W�CAf�A����O������;:;;1��ڐĕ��eM3�]�H禺$bT"vH-=?����^��I�H��%WP�����,H�7�%	��db#��� ޲���G��� F�000000000�����UB<v�����{屢�D1e����<x_�җ��� ===���טuM�i}Ur�}3!�����s��P�<� K�x$Ӂ%N��C��p��L��S��Z�Sx�6z^�;���� �8�G	u�Pё���z%��O�����O�h�ʄʕ�D�N����~��K�[ꓸ�&�﹪[�6a��Z�$c1���s����,�	8����P3��<>� �	����g�3������5+��~i=޽��&�����;8ji�� ���~�m��?�2�>��_��p��&��E1� �"3�T��4�����+Zl�FM"^f�\���{ܯ��jp�`�f�qK�hF�-�Km8,�W��OT��Wǚd��c��0�y����E�<����������A4�E�ڵ��������q�H&���Ll��l!�%6!O>�$���o���3	������݋p��mX���.l0��L'�P�?�f�@+Hpyjo�]�J������Lc��uY�+�+��b�����ӑ��T�N�\:/�kW7����x���8u!��x=���D�����L�����k=���C%Q���q5Y��xޘI���q���x��Eذԙpp��q3�<e8lղ�걷Wri���߶$ya�e��}D)�e��!��du�M�)��nM3~�J~�N]����������@2�p�֭X�f�͛��K�J92%�*�����׾�5���[3finR���3x��Tu&����A��z��X*�t�H5�"Q����{c����F33�B�^�bP���	�AM;������ Ӿ��Ű�)�0�}��S����b�_[c
7ol����ز���p'��m```````���a|���ņ���dR��ZY���'��SO=5cV$+��q�<�އV`��:ԥ��[O��!�u+nEӺ�l"��D�$(N� ۵}{~���,��dA��D��'�M4,�2��z�"/�:7�����F���ޯq�\�S��܍��?��|�;����ɄE��o]�+W4�+O��;&��6��������@��ʿ�˿`ӦM����Zt�A��l�o}�[�z&�x���=+��-��a�c�A����O��F<�A�տnѻ���O�t��u����i]��m_�h�΀z�C ՜�[F�]���E,�_t	z���e%j1o˧P��}H��#ę�i��6$�u^� {n��oZ�!afĕ���������Ϟ�`�x�00000000�a�޽������+Wb��c	�������x��Gq��a��oJ�p#uQ���9xk�0�j���i�G�h�%l�T�9��x�&�k0�]�E�K�&�N JuY4��$qx�,���%K����MG��;O7+'vZ�4��W�m�o�+ۏqZgI\�O�{b������2����e�4 sy�|���]w݅T*�K����\c�Νt��D_jl\V�����t1�x<��OQBz�j����煪�!<3ռ��|���;{���^)���>d��g ��j��u�ɳWG�x����s\������j��+'�XG'�ښ�a>]�������Ό������~ꕃx�X�l���&䋸�#r51�����������/~�
�7ոD`�`@�̎�����4C\F���BZӶc݇\3����E�,ڛ_ȩ�^����
[��ن�F׭���gȔg�>U�I���$���k2�i?�E�h�;��?ق��˻��耙\h```````��3�<C���vD�.scG�3$��?��%�h*a��/�޷��	���-n�\�X�R�t�`<U^Dx�o�6����5!�T��� �<��-���%����P�K@�b�j���u���Jsќ#�i�4%���:���:�4&��?ڌ������[�+m``````` �Xd<��ø�[<[�4Ye��6866v�*Y���w,�Cw-GKCR�G�,Y.�-�M�Ih,���eDP��V<I	�ony�<�^E�s�|K��M� �掑w��So��^��)�9f���4����~�s=�|�u��/��_6���q?{��&.�Ɏ��������Ló�>Kl̟?�D·�&���ٳx��/Y�k��;�Q�R�,��B0�,�c�D��X��.A6a2@*�q!����.sY{d��ל*�V:�G��(N�J(3���+��:��n�9�?�Pa/��SowX���5Դ�?^=��芁������A dB!��
M���l��������h�K�7m���]��w�##�����j���ۅ�A��H�X�n�D��w��ba���n�_�!W�=嗱}+ :;fN��z'P@a|�!�V\z�d*t17��h��6l��`�˽s�����w�1?y�ì\h``````` �������f�q`` �=��%�PSm�m1~��%��X ��W*'�9&����;�|��z�PM�����k!ۇ�44JA2�U����#ޞ�	�eX⍸Ymݜ�9���,��L�t!_oZ�b�&�]�=��|�9��f;�3+��?�i!n�&rE<�F�!����s�=��z�Q��q�ɓ'�}���^b���P�5�33���+���e�Ww��f���ؒ�Q���@<Yf�o����(FN�����@~����Z�$˼ͬ�}�+
��ۛ��ڥ7 ^� +���H���vxa��gw`b����BO쟝<K�m�+z<_�Sۺ��0$����������?�)>��O96����k��vї�Τbxߦy���]�e�k�f�P�'É��fq�I��0t�y$��QӶlB�<�
6ݎ��O��$b>A���0�S��>����p��ZH;�w��~�D����6��Cf�A	����s|!POVˀ�-q�W�1ĩ������ap4�_��F.o�s�����j�ʜ�8���+�d������uK�\[a��r�90��#��d���9A�9��MB�h��nd�o ��n4_�&�Ä<���c�/���aH7<ƣ䇖��<%��;�։3t�E�>����󮀕�	��b��>���ܮ7;�@-˛[\��6L�>�vQ>u�2���p?��i```````0�A��[o���@�	�۶m�h��nI5۸fU#%m4�;���8G����+r�/�NAin�uKoDM�*g�?�T�YJD�]�0|�e���IޖXa<�L<JA��q'�x�(_�%�`�<�r�gQ��F�ZV�u&n�Tu��G��;��#?�	7�={�NL�^l����p�}_~���}�̥]T�����rqu��d.i��}&�*l`0���/8�̙3t�ŭi|��Ÿ��V$��- Bv9.��&��Ro�4:<��1�$�wF��ݙTO:dt���3�r�DĀ�?3VW^��]L�M6��u��*;�"��{���ɆEv�ۨ*]��Rg��م*7qv'��+�v�������+����-8�;�o���������� :y^�d�%�����1>n�o�j�7�@��L:T�R�t��z������v�g+�����എ�ǥ��RK䢌�sT�%%����,�T���A�f#|�����&���3���?��y���w�=Wn�b��LE��o��C0/z)L%' ��>�e>N_�҅V��h�� 
tmmm Lt�*�0�ܕ�8�}�X,��b����>|��E)0��eM�eڛRe�-��y$����gF��5@!�6)g�30�O�η���E"ӊx�1{;���a��=3q�W�Fa|�*�����<W��J�pr�8{��wҗ����@�HgJ�ZҖ��7/�ɮQ�����CT �'����a��da��)��qgG	��#G.J���k��㊥��X.��H������pca��>	�W�<[�]��ӍH5����!Y� ��6j�L�s�V"+��.R;�R.���W�Aa�C�
>��] �X&v����('��� a��f�*H�}�\���lbomXր�nZ��=c8�9
���+�"�)�|:�x��2�R����Ű&+޹yn�؊X̒G-ʼ]��3W4�f�6K��n>?��AN�_���ԥq�ϴ8>��g�ʆŘ�<�� Y%�x� n��.��P2M&z�T�4��T^qzc�P��B�ũI�p��6:��{�C�<¡R�E���U
�X�!��J��K��Y"���x�=�Q��S�nB�).�]Δ��q�X���%����lO�e�<�g7v,�d�B�-�	���C�q	��K�sX�$[�����;��o���(��Af�&�/��z� Dz��k��=N�P5�������ٽ���%vu�-�)����z��i��C�y#��q	יn�l`0��������MY{s
�u��w��x�ͅ����̑BqR^�� Оju)h��G�m��&Ǆ,7�����C�~���.�$�4F*UA�ĸj���ɦ%��s��1z�ي���ta���U��8��M��g�7�~��4�s�nq>t���ʢ�g�d���WM��5�Lj��]�xLf-�3|z���s��#��Q�|�ϟ���\��z��N�p�����y���{�?��7(1%��L�Nr�'��p�6�~�Z�g'�iE����~�m�}�Mh��ًʁJPA=1$F�yH�q1�o���W1p�q䆻��t���!�)�	��m��d"�����m���=0�	�J���t�Ҫ~h+yGN�8q�WE5��������ߏ���߫j��F�,��裏��0�"DS��.�|+V���{����h�9��N��k��w.C1�(	��n$�>iu�������@�[�u'��d��w�u�o#e��X��o�$�T%DYU�+����lZ�����nٻп�1z�n�Er�]��0�iĴ�j7.?��>I'�;9�cfB�B<G}}=.5.%�7�{ ��p���KE�(6̲t�B!`F�yȈ�jҠ*�%�tsssE�J<b m���\%��e/�I�qז�ذ��W�=��2���b���c�9t27ά�x����ּ�]�/VNf1�y��;b-�0�Ϡvɻp�A~���xn�xo��\��)L���f�'u�yC+n�Ђξq����3	���X�l٤V?�K���R��*���8a��$'����8D�
]��wH%ڈD^����U��a�$������5�0�1�Oޱ�N"��v�F�9pR'̳��k���q����m-�o�#Դ�q]Ϲ�4��g�K�0]y�1j�Q��ݨi^��׿��3��c_p�l�����NR�F;W�O���J��ୋ��P?�tL���A�x��ߍ?��?�W\Qq�ݻw�/��/C'.�/��{�!ճ�-§?�ij1=z?�0.tϯ�/s�:�*����&�s�;�CT����`	4q}v�-��B̆�3�<����wUh�xr̻���wM=d4�n�-������"��M�p�+o���Em�DeA�$Xqjֱ�}_@��oc`��pȯ�3���\���yJ�P��R~��^ш׷�ɄF��9 ��hjj��2�IEzU+���M�XT{M1�(v�����=��3�U�֯_������vT�7lB�*m�9*a��	����30�˘6�Z��'߷�'x��;>	�(=�6�>'j�pJ�g�K��ꏣeӯS��(Щ�a8UzA�AE8H���3v`!zv}�e%ל�G��R�G�K��xGJ\������}�8~��B�T�H�&���+eCԲae�G]�0�i�����p��wcժUS���ɓx�p���I�'���gb+[���R�ڪ:}ai��Qȩ���R��쪄�(���~�R�)�wRO2�˴'Ӊi!��d��nY��F�DB\�QL0��
N���ˏ`�yoBb%�F�տ��+?�XM���BQ�#b�"������6Y���dؼ�>�����ŉ!u�gq�Kr����ϻr��]ߍ��\��rE��b�(P:�Y�a��(�!�����?�M�6�}�
#l�t�̙3�&�%��*����W=��6�o��a�L<ƧQ�a�����ꌊu��ת}��I�1�.��_�6o�<��r�>��������M��t4n��J�t�6���]���7n_��x6���4b�L��F̎f7��	�Z����l�<�u�If�UE��_C"�,o�Qސ˶�0���HI���%�%3�_}��zw=BW6tK	(�LOf���B#��b	�5v	��ṬX�?`�|yw�w/�K{�q���|��k��FLTϱ����)�,-_^��e0u��۟6rd�hU�KV�H����aVIۭ���Gv&S�
a�O��Uk׮�^Qt׆�J�"J�dp������L�*qa�����_�f/��@�q�<j��?��EW�K6,��d����D����{�a�k?r�g��,;_p��#�,2X���M�C��U� T
��HT��u���@DmЈ��F�D��c���}ǇT���r���]3+NW\L5�@f����Y@���]�R�=GP���߲\Y>ׯmƆe��00�|�(�3�$�b?T����(�ߨ�ՃNy�]��"Gb'#;*1�R?��3a�аΤ*/�uP�Ϩ��;��Ƥu깪��;^�v����=�eu�pb�4U������D���޳�n{�{��/f��v4��MW|��_I^n����б�� ��\��l��)ԯ��W|�Y6;⇜�RC T���#��WU�(e�/*Y|����g�0p�I�&��kP�Y���]�X�#�|�t�%Q��r�6AϞ�mߓ��߷��(�!��&K|o?<��ls�E\KKKUV.��� �;��Te�}<T�DR���q�N���B7"�#�S1���mQ�'�������u*m�"����~�0>����JT��P��>��3V��&L�9.q3����ޙ�zP^`�g;�N��r�[�6	�̎�!�-WM�?l�6�P?�d%�����6���!
�=4���{xY�,��g+�̂�м�>����� ~[|�4�b/�O�j,UV%�.#�!>�GN�b��J̫���3�W���������ܧ�e7���{��]!���z�	n����5s�@oذ������>�^|�E<��S���G5��EU�TϮx,L!S�;>ֳ��w`T#S�Xv��<�����J�O�|7�*�+�'K����x�{5��q��!ڄI��X�G�������{g�Ij1�ٍ��{oZ��}F����o+nEӺ�a�ki��$OR������P,L<C8䙳�e��D�nZ��7zy�"�^�0,�C�+�}�T�Nu�C:
��Itƺ�젅���k[0����Y��״���0��Ȟ̼�Dm�O��Mm8�5�|a�+�D}����-YG,��c�&m����C��醐eʗ�|uU�S��,r(�6'��A�,�{����'֑WD5*&�����b�=�3
Q���iu����_UáC�02Rݎ���.&dm�t�%�����c0�QUM��&����DP�,7�� �!>�d?O��ç^Gi��{ĵ�_$�<�e�~�{Q�x�S��'��g��;��GV7�rT�.�t�F4��9�Z1վ���t@�ߊ�#�/c�Q��:����6�~U,|��v��6���~.d
���K��F)SF|u"�|d��#'�諮�����ݍ�_Bc��t:��w�P/Ν;W��q�Xy��.ң011AI�O~��K�e�B��m�H��|t��c��_���n�[�g���@FNc*M%��R,TwDT7��kf/�J��]݄��Ҝ�:�7�D�iU:��,�xDYM�����ߖNPW�v7�@�kа��6X��z�����S�U�C��J��'^C���>���[�G�Oh���]	�}t��J$O��q�@�߼+W4`ټ��;n{t�3�\��_�:�Б�0�\�ǿO��l��cP=ttt�W��X/�9	��rsa����$<��˲B���6��f�x�g�ׄj���K�,��U�4�v�ߗ��aⱝ;w�s�\��G�/��p���4F�.L*�@��=��u�I�Ot��'a0�QU��k�!A�7��&��h��*�D�!#��05m�0r�M:�H��_~ڟ���~�{�'	�R����Yy�Q	eJ�n��n����VVݎ�ޣ�>_Ƒ�k��k����T�ϟ6ߍI%,ܾi�z���uJ3�����_�:�u
����h�!;W��1�H�� ���^H�U��X9��_���|>O���SX�P��QH>]XZv9�S���+��zn��ćB�}��&ѓ�Z9~�����̟�h�x.���k�َ��L*��5#牄�L[�8�]L {�y�D��|p��\���1^���k���5d��0«R �f��*��ey��n黨+�����o����]G��z��I��9i޿y~�Js��F���g���Q�^.{eqq8S�֗���r�!^ZYZ$��u;Ĳe���,C�Y��c)�oa#W�<gT#%������^t��EcGa��/��z�a0�Q5}��z,lM��C�X���*퉓�1�l��� �v��� �i�*�l_V��t�	+O<G]��z�m�0�'���ވ�s�1v~�o8�")ěYlF̛��D�sSЁ��t�������|�SS&߶m]�x* �*�që2ү���j�r�R�g�G&�WzX��"�վ�!U��b��pdm�����Ź��"���tCE�K(����U#�D}�I0�%�z��#��'�P�e�}�"�P0' {�=G@\��g�#�쩵�5�[Ɲ�R��2i��)C�PEt����,/�q]}��y��͘p'�	��s
�^�vѵ�� Cn�����5��2�8�[ӌ��wa6����x��g���4�|�r�d��jΐ?�<^y�I�{�F�>�P��a�E1�l۠
�4a�/S� ��,{d�X�]Q��Hs�w����$���t� �FidD�9����k��L��!}�!*�8���Ô�2�)�de�񞣠Kº�Rp�t�n>��@�W*S�0�31LG�u���F�RzE�
�U�Œi�-��g�ӕ��2�G�E��k����t���{�7��X���[g=��~���'2�(��#�������.L������/��^V
R�d2Y���;.>�a�����ҋ����"Ųz�B�:�QD��������)Z[[QM������((I�e�M�����3��c�rT�@7�&�za-]�Ё�3_̈́Y�:m¶���	dWJ�c���3���@�C�nKK��y%�V�%����GQ�e�9�C���1��G���d� �PX*0��`�3r��v�B�-�<Y������w�8!WLɪ�[�LM����Q�6Ȫ��o2hhh��u�"+e��(W�n�<�#�*;�jׁ/CF�E�2�Y5Z�S�e$ZG���Mp��b���Ums����O?�֙��;�]~������T�@�^T��L�AK�ML.J��R�S�"Yߎ��c�! &}{j�ͱ���\�����,��y�P5 ���G�A�pGQt^W�08*t��g��<��q&���G��oa~��y���>��}�ل�8t�Ē�4�5&�=8�WaR�4\���0Y|�<š���@H��ջ����Q��2����qda"T�"��8�D�wN����;4eX�mձ�2��b�f�3lDU���uH%c([��C��9&��n����.;ݴ�#H�� Y��	A8�8�N���� 5-B�v"�b���~����֩��(�2B.�+
��E��*_��'Q��᷄����Ѽ�^ԯ����׍L=�;'O"۵����+P�`	�1�aò���s��W�0���I&P�b򿺏��C9u,.;�����"N��S�r2I��*�,�F��tߛ�
5��<s��
�sȟ�j�=���dq��S��^T�L Jw��m&j�����~���BM�Z�D4Q����y��rC穇pYQ�g@~b	ꓘ�� BV5VQ	�9�ʞYg���0�l�	�W����tyo2����V�`_�����M�����(�&G���1�s}'�맶�n��u!n��/�;Z5��#
���PuNe�T�c�!l�b�����|NCT�:u
[�n����.�HB¦�@8�<_%dBN�Q�J:�Q̣tD[�G��v���̌�b>?2s$h�f=�B�W-���c��Cm8�54���C2GHQF�YYԃz��O�T�yI���8���k!^Ӏ��Mԫ��a�#�Ե�FJ���GQ��p�p\�Y��N��M��c��+�5�l<��P��"k�d♃yJq\�M�{#���	)͢Z���%U��QL�t۪�Q��x���'?����m����_Ǟ={�V�g�#oi�MWd�y������2�S����J�rX>�q�T�HW��e�������L�S�ڛk���Sr�/<�7�١��0N�{I�Qep�H6d"b�}���RD��)��'*	��)��L	�)�DQ&��!F&������f�biV�7�pR�8��I��ҒbW-��zx�#�h�L�l�D��S��ŔA�>��,�,�'*jkk��m�B�D��r�	 �d�HL�M�e��j�U#ZQF3UeEAT��@��@VͦV����=��g�@�)�-)�S�ǊOY��Y���Ҁ�$�^6"�=�$1�`�v��U�X��J�udC�TB�sU�D�$���qWIV�MnGGhB�CBǇKP�t^�zd�./�8D��adt�C��)�*� #�a�����_nЩ�"�_�jAT�Æ�e{�B�n�аK����1����Kݳ:�@K^R��zL�@/jM�	���q_[�'��ߒ7ጽ{ޒ+.!f�fa�q`��p+�B�i9]�Zgb�ǯ*��"�y�����ʔ�%�ե��c!ٸ�z�(N�+�v^'�9^�P�#����y�5���7�����r"�a��à������U�������AT��m����F�e�g�+<!��wF�fDҍb��!ٷ$�XO+T�*Ux:��u�,Ŷ��Ɣ	t[�Mf�'.;�X1�ōvX��X*�;�9d`��M���C��%{ѣ�S���SӢ �t�@Y=eu�5���%�%�tYt�a����7�σ��0*at�L�|�;��5s�@3D����}�ŏ�*���W:���E�?g!��ˆ�U�Մ�Q��$����Ӳ8���t�0ݶ�d$(�s�<O2�\R����jL�@7�%��W����h[��K.Ms^H+и{�����جxɆN�"*�"�氡,Y#�
��Ol���'�WAv�ɆŰl�u^�e��sy�ݿ��ڱ�/S7����0�)���=�=�3*�I<�R�e� ,_]�|&;B4�!S�u�Z��o�H8�K=�P��1��#~��<�mջ�K��n{�!>�����ti��;!vHe��`�c���>I�]����f�UH4<�����B�=���<s���KP�4\�aÍ7՗^�����ʈ��1��^Q���m6�f��uXx{g���䅰-�^9!����NX�>F���]�H6�0���ЩiaϢ��R�dC,�iT��:�Q�K(#|ݦ��Y��3�ʋ@����Y�N|�eD�Z�,gU'��3�՘2��O��Y��������&�=^�F 9�w�����&�q�:Y�Uf~!��eeF1���Uk�T�L�XM=�fN"p-�e��<OW	n�A �d�>S��D�L�#�3�æR�eq�m��퇕�ᐑx"A��q�nM�t�M�,U�t����E�^����>z�(��ƪ�~��.��A�\����=;2����X�Y���c�,�&��gZk�����>[�@��FS��d���X�t�r��m�a�|�>Kǧ�GM��<��2B,G�_���<�_ⱄ�vf��vv|]
��~F�pSqf���u�7��s�@��X�����L�����U�3ϧaa�N&����;�;"�Q�^�����&+�u�f)ѵ�b��vd�"�<?���#�ϣ����ĴC���~v���X�y���`�a�:�C�����/)S�ƈ6�Kq�~y��ny��
x�БNUC��F�u�*R�J/�(娔L�ݛ�@,��cv���#��r��)��8�v�ŧ+���1��M�1fRS���LA��J<ƎG9/��z?�@T�D2OW�2�SR��D{�@e�!׍\LF�>�<��,.;Ȉ*{���a�%M\`V=�zL�@3nl����/������Q����Q7_�E���*[0����Wŭ�P�H<6��K�/S����ޱ8�����8N8��La��d���r���� 7*�L ۟�Йo���+g2���GQ�U�2��B膔E���S��TF�ee���,�d�{݈�ʄ�rjkB�W+B�鬃��Z�f=�L�}��#3ݸdqq,W�d��5�̃'؀g$��;|�G��S�Tk>��Ojt�e�d���]<G��_,B�%婴Х/Y>���i�՝U�r��'{�TC�3�t����Bܗ�3�H���b��5����
aI������վ�2QT�d$~�h�wC52�1�}�d��eA���V빑�b�4p�2�.���b�m�[��͓���,��|�9 p�;��aLܥ�5J^1R-�`��TeTB~u�.O]}"�{�
�W��W�E�[\n;�ޥ��uƜ��9�I�X?�Ȏ���F�t�u�B�I4�$dꮌ�N��)#� ��� Ȟw�ȕnGa��ژȐ=����z���T�Ȳ���K�!�sS&Ѕ�KvA.�B1�Ձ�ܜ>mY~�pϻY����`)?$3n�hd���qԏ����Ht%
����l�6����(pSj����k_���9ŗ�+νVD��N湺P� �c"	�d�De֤4;
9n��"!���IPW߂k�u�kG'��ΖX/��4.g��kٷA$�*�-�Qf�&Pu� �U�(s��K�5�1�2������sf�n��E�@|��C�݆���(L!����U�ta�@g�S�'��dy1?�R��
(\���e�a�zy�[3r��&
��	�J	��.Z��l�w��GECC&��Ǐ���s2�v�J�Ʀv����baj�m�(��k�O����p�7��k��Z��y�����Ç��7J�-��(e�D���nB<^�I�{������U'p��0�e\v�2�Ύ�Q�cf�Tg&1{�<w�y�y�N이�� ��p�Q���C(յ�"�.�*d=�j��XI#9��T����� J�	����xef�l[�`8	Ɏ�-S��_>�rQRy͇��!�ɑδ�m���cbb�q�uQ��� ���c���X�:i_��$s�a�}��=�ӧOO*+GMm+b�y�p�	;�o���� ��y�����ݪ�Y(���/������:�X6�#���:�b�g?�Y,^���������b�֭��&���Q[KF�]�!埗rEXB���}��`�d�2Q+J�3!1��2���R��e˲����N��ϛO�K��h&Q��b�lR���ѩʺ}�=~d�ZV�0sY�U�*�l�kU*���md=��ut�ݗ�wS6� (���pvnh�P�*|&Ce.�:�(�C�i_��� ���aP9.\���ݏW,s'O��H�wb��N�@3�Ͻ�A�b���N�����U��k6���d��-�o��ܣ�CgÆX�f͔�X����i�{�ӸjMS�~m1���}�:*N��:m�kK�N��t]-��#Py���L���y�>)�x��,�n�\R�A�e�������Q�@n�\Y]���,�寤q�l�&#�*5[������F{�>Q����k��7�8���X�+.J~��'� ^N�=s*������0;J��^�8�H���L�D����غFK^e$u�%��T�*g2u��P�6*�,���}���b^��x��(��L6]w�/[2%M�ܦk�d��u��߃tr����`�� �x�+0���r�7�C�P�L2|���9?��+{+�P1�����v ��݃�����J�,�����9)C5��j(OF��ʞ<�R�is� �P�پ@����Pi�O�Uho&B�4����Q���V�s�L:�U�H�a�&"jS��3�fE�����3����'T߇0�:���u���]���$k�Tq�≚@9�΅�{?�z64�a�w���&�{��S뱹!"�eL�@�N O&��tH�g̖#'����v|D����h��'�D���?�2r5ɔ��'�D%�a�T�x<*U,e�n��$�9~2�@�#e�+�J�	1�����H�p����~����>X��H&;}��_U*�:�%���}]<Y��CE���0W��ȣl�R>�kR�h��'/�
���H��`W�cT�g� �%a�V�gGwߣ>#�S&��6�&
�����i�?=���a�$��]~
A�ZP��(d{���d}{����7�c��~����ś�*.�'F�:O;�x����64�l�a$Y�~���MVa�?����.Y��7oF*�R�Q�Q�}�����WT%�`ꨄ�L�}������s��M'N��L@%b��8��#��l�¢֣_�K���v��橔��_���S&Н���1ڵ�%.�,��:d�r2'G�q	�܀�����jm�7���#9�:r��a��,%�.�V+t�
���p ���JUK6�o�z�<T��}�t/W%*��T���������;O!��j�.�bwJ�{���蹷�=���A.�X/o�n_Gvb�x���Tܙ�3�&{^�΃Qm��Q>L��Z����җ��Xljk�N��d0�\����}T�CamM�2f�s�=��lg��]���)��l��q�@�ʀ�Y�h8v<݂��D��#Q�f��� ֯|�7ޏ���a��36�v�jF�]"M@��u��ܦl�Td���_q[��\G%*2��Au��c��Q/>y�G
bH5-E�!�`b��,�p�R@��;��A�����oS��/�������.Į��z|��E[[۔�!�饗^�SO=���~��>��Q�����Ƀ��ݵk������ѣGq���]�n3陎
Ug�Rb��V��K�mY}d�L%#BQ:U��\�kP-�7?d�1���2�&�ə�,��mB�u��=��<�<ӊ��@���H�9�>�d;�D,Y�y6�KdZл��(�r,δ���b��J��ŭH��*�i,d=ya�bY�d:�:A&[f/@al�?0�H5/Ǣ��_�D�h���oZj�\�D};��#�_�hE;����}�g:���p�WRS���\�cǎy��f
TdV����E���������_��W��pq�v��ߙ��g�tT�����K��:Rz)�7�7�7oޔ=��ԩI�%�=�#?�w�t �+�ُ��)�q�s��H�N:�u乧�d�5 �/��W=H�T�/�M�Z6}��0t�E��\��en�����ݨ[vSY�FA�{,+_q<�-StqDT�p��<�sy��'���2��,����I�
u}i��qZ���='�3�spl������M��*Qp��$�����Fh�8�v�]~%C��r�̇{jP��Q�F	�U�I���E+W���T�޽�*�L�-���~�'�xb��'���AU��C���ZI�l!ոM�?DMDH?�6ik��0rvJYס9O�b�#�9��M�o�C�-e�b�!�Jd�Q��uiduѥ	�3�Ϟۅ�p'����а��H�o�t��v�5�]ru!X �5�:�Fc��!���T�򑺘ЩȪg/�J �.3}���@��!{�'�j��ӱ/��xW/u'ڌ�DEU����tҘ�����~,A'��[O�^T�MHwz�z��~Cb6PB�0��ޣ��;�T��PK$ �����|:a�œ)|b\U�z��$a��.�v�E!;�����J7��~Pz�z��%��j�z�����OO����� ���V��[M���	�X��=_F��!���4��������y2[tY���T�72�q��,FFF��~	������:zƱ�-b6T�����4��G����[��3���g��#7�i�mH5��ˍI2�$��� ���L���#�v�Q�Y'��|�0zv&�O읝���cv�䊲��un����i@p"�Ǒ/=/�(�d]�G�A��T�(�}�U��㕒������Z�����?L]�U�o����#�wJ%�q}�Q444��طo��50�˨
�&�u�׮n�	�k̑]��y&3�=f$~�����sgg�Q>c��̣~�-tB\�����m�iņo*
��\��s��_�B���ޢ6�\)��s��Щ�<��!F�c< �|�m��0�AT��'O҉&Sq�5�jN�=��w݈K#�Wu��011/�K�\.�ӧOӿj����W�����k��#j'Ṽ�~�ߤ*���AuQ5��p?>y�Rdj\O���R��b�Y	O5,�"���!����ζ��p�|���B	�n[�F���23�ݚ�GXEO�O�����7���2�����e���ݱI�k����R!� ���B�]~��*Ŏ;�D�j���<���t!JÞG�3���҉#7�4�*s&~�?.�V�S�:����`��~�� Gsh�M��q;L���������+G�K�:U>�U�x�1Ā�q�*���]�5�(�SlD���۪8�42S��� ��dq�u9�]�&����Ʒ��ȴ_:����s:5^<_�>}!�㝣�� C����eب����H/�!�'Y�P�?�++/��f`p�C'�Ȉ�x\�S�0*j``�����<vĢ��1&v:�牾6a;AW�)����3�>�)�.Y�8q{�`��/�lX�x�1�O91/��揫��JP�FLL�ʓ���Os��^����\��^�o���H��@W��W�,^�c�!����==(	�i�`�<t�2b<Ug�?.+�|��t�G��G�0����3+�a``P}T�@<��w^7�q@ο��QD�nE[�j׬R�Xx17����S{^Vp�NZ,N�P�Hz��ۨ���S����T�B7�6��du/;^,`��~�|ٽfB#��l�V�A=k��Tdk��0�7������(q&�4�3:�� ���F�d�N��];��Co0�!~d�Tm��L�œ�e``0}�*�~�@�Grh'������%+
��|���hX�^�\��7$.Y@��[]�o�-�x��t2aM뚲�UbBQ)TdEe�Vi~a��������t�m?�@s�/6������#�vbY����_�"&�O�%��{�������0��'ap����Ig�W��!�I����R�T��,�!�����RO�3zL�J�/L`ۡ~�s�/̣l�Ǒ���{�(���S��s���č�u�?E'�z�<�Iebg�͐}�9�n����m"�Z�jD�n��7C�"����l�tʶLu�������R������&����`b!�ܩ����B�Bf��HԶQ"�]��A?]y����ݎR~�ˇ�����1:~y��v<��s8r�]���ď��.S��+�t�\� �,�~)1����2�J�	~�Z'>���v�Ů-��;1p}{�l�^��]a�y�%�(�Ǒ�6����d8i��1Ź�m�p�n��B��6����^����b<Y�,�L֥�ٻ���v�g�۝�_�ɔV˛oX�my�6��h���"�����3M41� ���Tu�.�$t����F�`��L�����_�H�Rhmmť�Y��`����������`.��z��~�<?�Uk}e����u/�g�D��-�Ru�5�T�@�;���C$�t�_�7`�Y�s�,�
�����mE���b�$���Qm��c�g�2-�b!G;"�����Sndd��h!����6Ƚ����;$�n�ca��ky�� �v�����7�����������@�������G}d�#n�3�:GUS�A����D �d�O�l�.�����)5�]�V���C� ��\)�Te�DJY�@��<ƻ�oϏ��E�<�Y�2�@�60v%�E>?�%�o��c���3����������@�	4��o��o}`��q�Xp<Q�u�Y��g��7Y�A�Az����v�f�D��:D5ᠹ�̜�ŋ2AK#����BϮ�Rf�͟�vC�_��w#�:=�5���΍b��L��l``````070-��g[w]��m�Rr	���zF�*�.�h�K�-Ւ�6n˱����2�Q���H����C<ВC��|y�Ҋq=�Mȳ�1���Md;�x&/BM�]X�{��%vOi�L��������m���?���i!�d2ُ~�A'6d<�`��A�hy��o�Lc�����#����Xt����<� W��&��H�Ώ�Q�@tqĸ^��<F;v���`�Y`���%^K�r�XT�uJ�H��}g�����s�B����<��޺ءm�y�C�k	tN�v̶�O �@+�(Q?ƽ;�C]�5o| �T�����M�V:�Z��Jy�x�{���s�Wg��g�9GT��e����I���<h``````0�0-����?|�wmiG}:�@�;���E׌�3������x�pf����l�9�ȏv���@ڮ��eNv����6:
Ig -{v~�'~ew |#qob�WJ�o��RĚ)�ey����F���5>F���@K�
M<4���-�����;;?n�Ar�s�ό7��n����ȓ3� ���O�����h���h\��9Tb���[X����X�Եg�#�M]Ąy4�\�r;g���w����H�c�$��7��	�E�>�1L�&���;���棽��#l��:��z|�	O�x��^���6E�m��r�xG�z�>�Z��mԴ�U�fT⅃�l�CUޢ/�	�~}���/ӕ��#�w-�w؆׵��K����<=�_�����Q����@bw�|��,���VM6໪�I��?�P �,��|�h~�`_�����B�O����{и�N�\��H6�ː�V��N��#��7?ڃ����K��;�9�+��E�R҈�W�-n[�<
E���s8tvDU������,Æ�}hF�Vj`p��{�n<��ct�i%�C�<�s�y�wS�Y�艝�lj�����)��������.��Q�����[,Е����<�����i�GPӶ��>n'�i�F��YU��b.ł3�q�4��>o��9J�D���!�xyy�-�:)��kL8 �j�<��%��p�A�-�{z��^�y����`aݺu��g?�իW��`�����>�y晋C�	�vg��gO�o~g��qW5Up�|;h� xq]��gX�Hk�Z
��{���-�����0�'����L���_�^�.��L�ͣ�tAF��l��UfT�.�P��q���6q=�6]6;��9?�������4a�|K`�]0�aYɼ�����tN��;q�ss21���6�l>_^%��O�QV�տ�:O&�X������:/�k��nQ���|*����S��E!�d��]G�������Y�D�Q�rk]�+R7ry�h��ע���� �W�}�b�.g=ڱ��\��4�dz#2��Ez�z$�P?�V,�(�.��M���Œ�.��,�R*L�0�K���؅l�>�R������b7�]��u�x�	�w�x;iw��ʔԁ�Wr���_�ĶC�(a````0!��S�<!�FE|D�
����;��/>�(D�����'�L��b]u�T,_V�J���z����ux&S7Y��ԙ�;��B�	:����W:pՊ\m�.�$>Oj�\u�;�j��H�-V��c���#���ȩ7h������#�`wjې���x����)/�e�ꂝ.��^?�6i�8�\�i���h��"��.�é�Crŋ!�@%vr��h\�#D�w�I���]����]T�60000����h���j4��7\GJeu��/#k22�"\:5ZU�N��EQ|u�3La�����ʑ]�y����^ש����p������p�4��3��ދg��\�y� )�	������O�};^���ό�g�����="->8��+��"��g���!&��nP1���[��B Z���·����]̄W�Y<�
K�m�
[���;���v{O�����`�B����A>M�|e$:�JV�Nm	9�b�"��u�(��<ea�t\dy��Y�T�1���{%^K1\���]7Ub\U�T��zl��W��b��N����.M�gd�簔�Y�8K�W�2%WpV�m��X��L���1� &�J�C��9����&�Jtਥ��R�v�!�%��,^����W�c�z�Ӭ�1j;M�~X���+	g����� �ge�p{Nd�ot�Ƀd�v���©"aa�	�0>?�*�#~|~"�(dU�Z�^�e�uՑܰ렫���vU���)����Ȼ��bXXy����"�����r<��9,����ڐJĜʁS�=�Wԓ-FS]k��E�y��m�S��"�h3j^�d�"jnQ��x�1��ن���ȏt�ju�jeҬ ��5d/�3��N2@y�ۊ� ղ
��7#C�\�Юs�&΃v�c���]8h��B��v#H�)�/�c�ՙ��%J�Y���^�;<O�y}��糁���\���p*¤S8�҆)�Qȹ����Ĩu��Q��*UX<O�U���ߨ*��|d�"�-S)�b<���҄��ЕVW�>�E'���/�ł�j�	�$�w��V)!��
25��W��z4_� ��W"�Hy���_M�:ԯ�CG���c�P&�1BM�/N�qDU #�NU74���o%jQ��&4_�1�筣�����+oà]�OR�j�LV5�A	��wW����n�|������;��g�0x�*�⨆�UdQD����0*a��%�D!�Z����4�:���Tsq���UJt�����3�y
{N�륻���@���C��D�C+��=�_iU}A��Oly��9FD_�G��-h����i]$��E�'k�x���\�{��ȏ���ْ:��%�`�|�ٛ��~=iX�a�ֹn�Mh��SH6-1��1�h��È�u���G=w����b���:^-J��I`ה\��]Y�о?o胁����AD��T�ix�*���X��>"dDKW7>�J��R�u�6�NGu�M�wXgA�.��+^�篗��GU���r�4�q�\1_�~ʞ�KB�	�B[w]@[c�|�R,hI{�J�E�O�)<ȑ��A��&��i�]6y^+�`'��IGݲw!7p
=o=JW�ʡe�<sA"�/f��@���L"�I�T߫3�p*�jZ���"ٸ��[|(���P�M�w~
�b�G�yX���s���u��?�7��܁�vu#g�\��H9���(f �_1�H�Tq�1��M&��S����:��c2�L�t�(�s��q���G���4V�\�x<��[T�uDYv.�<�uSuH����\2M�;��c��GSm�߲m����-��< ����>E�kQ3o=Uu�#Qs��LM#&�M9�/�#�|� 1ee��ryS��nٻ�jYA���u���I��Kn���W�:[�
�M��q��lj��`�ݶ��P?{���<���������AE�	T
���.����lccctU7��ŐL&�_}}=��܌��6�R))�����J#_�J��ME�e����)+�ߗ�Ӳ:���������{��X�/A��_��_���Ay�����`G��U��by�{"�h���1��Ԧ���h�K����-Ay�l�皖UHԶH{Z�^+1� ����qn���q`U(W��]�L�r�?ɱ��g	�,�x��@��Ay�ć��9Y7�����7��X�`�<y&������=�߳������03
���r9ttt��w���Çq��)tuuQ=::J������@���c��唠�]��n�8����*S\EE���C�Ї��|~:5��ʔ�0r�:���kx饗�zӦM�>����a����gB�U�VH����3��Wf�����h��G�ݭ�Q�����G]Ʃg��n�L:�I�1F"U�X��S�e=d�E��$6ٰ����Kf�w�� �w�(	ۖ���^�!unL�rT��i�d-6��@y�z�J�� ǆ��<��ӴSc````` "L1e ������u�V�رG���yppPI�T &D�^�x1V�X�+���]w�lق%K�DR-u$_E���tR�;�H�F�y�H�L�U�ɮC%Ϗ������q��i|ҁ��w��D"!���
�g�����]'չ���p����IJ��It}��mq�ǖ늍�j8j/|B���(��/��+�i9�O�8r �젺[�	�G\9B.�ˢufŖ��d(��y�݇#P�����2���DO�ىo���<h`````P	xBCҏ~�#<��3�4uwwO��
�Z����z��r�B?��C���?�L&C�EQ�e�5
9�AG��:�ȟ� �}]FE�UJv��L�z��:w�^|�E�۷O�hr����d�"�a|P�^U�C�	����=uE��w_ߎ�t<(�Z�#��MX�bn���ˮ�T�#���C!����IЊ8e�Z����Ƈ�:�+{?�y�_��06��_#��@U,�I�x�����l=��y60000���<%�����L��;;;��b
@H1	!e��C��F�������VN�I��VXGVv����+Ckk+%���TB�Ŏ��N�9�:/,�j�BVO���1�4��s���'OP/ܲ��Vȯ���]��X6|R�e�8KW��#I�N�Q�uB�G0DRL�D�м��@Z�F�x�B�c��?��«O�+������B�}'4WTP�]՚���ֳ����ntP:b��ꫯ�����}�vj�dr����D�I:B���Ml�+���۩�u;�*G�RIeDX'���Q&�)��.O�ɗ#^�?��?C����G�Ĳ�������+>��k���P�}�h�S]Y|�?Ob`8�߹k9�j���;i_}v.D���F�P�pS�W*L {~/%�t�LV$\�5��v���������~�^�#�C��y�zuK߅xk��<�a��_��.��/|^b�� �p���	�����Q<�z'��a`````<� 6�d�����@�J29��o�>�j����B�4�}%i��L�u�io��&^y��8G1;`�")
�a�)�bQl�UMU?��R���X~%^WW�T^s�5�|T�3L�VAwmt*;�׺|t⤘FoFh����xd�t��?����M��G�= ����#>��H<U�P*�8��w~B�8���d�{�����-~-��l��-q1�TLI��kǻb��HԶ"V�$�{/F���#8�%�����\��;���:�M�����م�1}Cg````` ��U����ϱk�.�AB�o��6|�3����_O'����aY!q��.��n۶m��w���_]J�e�		WՇ�'~�ل5>����D	'eu���6`���%6�'N��&+d�����')骩�����bѢEX�t)֬YC]�����e�9���	�&e�RG$���u!��	�$>iP�a��\'�L���s �iT��{���@��_�i�LP%6�^� iH~�����F�HO�щ3�Y���ވ�����*�"��J�����"�H��ʏڤ�MZ!�Du�z�_<���d�Sy��ɼ���K�D>^���|sV�����JԠy��R�v�<�]8������g��lQfW����'����(v���De3����겢:wW�����$ �QDap 
�<Q����ǋFM&Kbd=׊ƅ+�&!Q���`�D��	85�Q&hhhz��������v�N�s���{������T��Ug��;��
�B��d�ݷ�����f$>�|�;���p9�%{R��%9��0���C-����^_����[o��D�W$�X�< ��x�b��G?
o|���Hx1��G?�Q9kx����'�z׻J�k���p���7����/�fCB�����U��	�0;U��=�y��y�k\�'r8��׾����pF���˿,���&�v$����g˺ƀ���?�#�k���6�m��w�+.���y��_��O����6����6̇����^�WDCn�3�������>���EC|��b{ٶ�u���x�e��y��^��c������)�أi�@�w�=���ο>��#�����x��2�i��[��3w\��~ v?��rq��ԞX8�n�}W��;���{b���=I���*S��m����Z�DO(���>���b���=��yg��}�83H���m�.;k~{��+*�)]Gک]l���g�����n���u�B�P(Jp�!AjR���7�_��_�$�*y��cN���b��ֽ��/�k���$�t>h��dl�ҥ��y�`�ډ�����-I9�FŔ*�H`-!������?�AI�چ'X`��o�[��GqDI�0��+�H�q�e$���K@���7��<�H���+����r�trhON��	��o�=c�@�c�a�Ŏ��Ā!$�6|p�s�m���ЇK/����Å�vޱ�����S.ƀ3���~N�<�F �{h�8�w��N9 ����9�W>^��wl�����Z�F�r�3��ZQ|�q�e�C/7*袖�r�T�5$�]��'��h�P�&�	�m�M���%���[`��=a�������o]�0�ض��9d�Ά	�`պ���&����r�VP�P(�.�J�UW]���������REF2-�s�byQ�~�s�[��}tʳ�kz$wH^�>��R�D"�^@}A��.�6��P���?��rd��@��;��;%A�袋D[Hj��	'�P�X\/��Y�<#PI����݀��ֳ�1����������<R
��o}������G���{�v��/|a��S"n1��]�~|��-��]��8�9{��P��pQ�b��8A:q���k'��0�!���ӆ�;�?���HIE�`�vز��r�n�g�R�u��@����W���s�6��
�B��� #K�+$���{5�"�M�/�m��! ������sJ����}����.��Ga�_B�a�Z���mT�i~���P��/��T�%���~��K�U���B6�>ǀ�2��rJ�A��� 5�E���튝(������-[V�f|�Cr�B��Y�9�ca%����Ke]��h$�7�v������N;����a���a�LP-�b�m����A�*�u�B@U��k?��\��,�h�d�*L�LG�-V�)P��Q.ōK�_|�2xJ��V(
ŀ��:ܗ�\����%���U�ErN��U=���,Tg����:�t�I𒗼�T�<�@�Xb�cT:��a7�.�篶x�'�Ehp����s�1�׽.��1/v
�>���˴m�L�!���`x���lۮ4-��m�1��@�c�cy?���BX,Py��A�H�1^ J�Xy���N�4;߈Ux$��X��,Mxz�8����;V�Y�9^|�"X0w&̜�#νi{�ZP���[��Y��-Ux�\Ԗ>�~ ����[4(j���VR,�iɡ['+4�	{90���^��g�Uo���:+
�b`�	�y�dz�UŘZ��>�믿>N�U��s�!�6�N��	9���#�yp�ÙGN>�䲃�vx�	~b�,�T���f�t|8��b�7Χ���WT�_��ז��PI�����o~��٥*>�o`�HH��0Zŵk����m��W�҅�`��V�"��
3���$;.�Vd$�p �W\Q�r���c���C$��؎S��pX�-�F���g�����^�7�y�~p�>��+Π��2�~@]�HW������~[\I6�� ��dbM�6>fڄ����".�u�|l��z&�3��x���On~�l�{�
�B�Pt%Uwۤ���m|q�|���O��%a삷��me~�/�{���
������R5�AsH�1f����1��\�XjㄑlrX?�|��I��آ��1�1"����9��g$먼b(����D�>ӰT��pJ�t��b�����Z/��&���h�m����)�$|�K_*c˹��q��6D���|��[cM�-p���w�oV�'��|�^p�≋v�,�iB6�܂DEX��eݒQ�ӧb�=bn��HyA�����&�a|�6s��9Q�1L��hk�����'6�Ony��������B�P(�E�xV����.�m�c��s�=���Ȫd#6@�1�%������:�Z�z�ꒈ����/J3YX y�~�O����N+�ѓTh̃��8���Bc^$�8�vl�6C�����:�V�A��6b3��6����]w]�!����,+�&[�����hH@�8`ۂO�G1-����>������N<jx��`�]0Fڇ= ��rVa��� '�w�|.��KqL9�#ȡ@�;�m���y�q^�nK�b�w<W޸���N�P(�a�	�ZU�X</�
�FD[��mUh�'I��l��D�A�XZ$p�S����"�]`���T^q�;4(C��c�9��v�g��-V/T����⏻��/�fa��� ��#���_�b;�m��Xq��:B��`gU���0�4������?��pů�+�]��;���}�>{̃9��(�u��B�85�G���|�-TJ6Hȸ�N���+����ݤlٶ���N��ݱ���)X�B~m�P(
�0@gC�U��@ƀa
4$��$�6�#R�1�����/?c�nW�f(�O��f}�f�@"�����n�G̃�
8@Q.��
��-��1���mmHo�7����`��/�c�'��_�1�8e�w�7�p����o�"�2���z,�0�.���p��{�IG?�ox���`���|�5HE`	]��^$���W�󊱡����s8�	��ӟ����-�ȓˎ�/�Z	���xf�`/V�B�P(r@_�r�"Ш�a\.���P�DQ��	)�z��S4M�'�Gu�_�B��]j*�H�P��� TA1��%�tK1�hg�@���pz�����e\7*��!�a�7��Ǘ5��ڢK�3͗:��@�T���{��Bc��\P�����X�4��8���Ӗ@S�X��X����p��Ň����k>�_�i\��p� ��R;�L!GQ)܅evq�4t��4�E�u[o�eOo*����%���{��+�7
�B��*P�j��ƀ�o�
੧�PC����H$1ng�h�OW��"�|��w�w�\�1��>�YB0�z�}�)?��8�NU�Z�Z
'�ې�"�ö�Th���$�^��E_���@JImD��Uhn�1˨4c(���t�Me^\�Q��YC�y��}� �[��֔8S�s��:p!�O��g�����fCu����~.�������t�._;��*ԅ��c���"1+Vm��Wn*�������&��ݏ�+�3W(
�b��	�b$��� �2�������{�O$�n�Kcn���bm���Qݍ�g���ս�-o)I.�G�x`;�/�T�����d06��t\���l)�~xI>��4R�z�Y8x���Ou�R3s �<��6DR�1&�����i�m
��`�J�}Z"l�����M��.��ΞQ�ځ-�ҋw�;�7��mN9q��Y0g��{Y�q��#���4p����!+�n)9yb�8��8�'6��1�Y�P(�Q'8P��|'��?�C4.t���	�o��]�[RX��Ŀ�͛c�����1-N���}�$j����I�v>p:<$Ѹr��nG��h�]1t�'�-�r�f$I�kLz9�k�c�o&l�!����#v�g�q�8��߄�9�	�c�Q}��x�.;-��ؼuG_�$�H��^4�$Ћ&��]g���Ο	�̝U*�H�1��|�b�ڴ6o�u��Sέݰ�Y?A�'�3.��	=�e�f�B�P�6x\,*��{��ʁt��<W@�O�%������wK	RW-�ض>|�icT�c��`Z�$���������G)���C҈�φ'p�ꌪk,T��~ӛ�$.\��	����ijz��q̸H����|��agUh��YZ�W��?	H��m
W�S>(����ѧ6�ؖ�&��.�f���3a���0{�4�A=Ô1��Ψ o����?\�U��J�
�B1���P��U�O|���?����T�1�HZ9䐒H�`7$rJ�v��N�E1��׏��|6���1�8�a88҆i��8#	]T�c+	�Su�?$�88��B�q�.��S�!Y����sKo;V]��_��_����d�cm ��.�͌�BDPE>��3K���{Onc�s�J�3��h�[@�P(��\]D����?��ϕ*b���+v���/^\��p$�6�CR���>uUK�b��;���ɘ؁@�"�Ƽ8��������Mu�8�?���;&��w�}�o}�[a1���� '�vPe
8�v.06	7� ��`G ��S����'��"�����̛�U�y��Sa!u�4Z�P(
EgH���]2��_�rI蚖�F��8��_,�U��=����}-�ۿ�[9��������/��0�;hg���6������g��ÎKiD�g\�ERY��/����1^I0�N�'c�����M�a��)�G������8pV��w
���1���_��Z�P(
ER	�耱������K�S�xZ��G�N�S{���W�We�J�n��.�́�kc;-]�4�K��bqi=��t���R�-pq�w��e���v[2-ō[ !��In����C�����؀B�'*�80À����A��o��c��X(�V(
�B��PQ�D�j1�����p�c/�-^�|Ŏ��1V	*�{�w�
����`��O��z����_l9mU�0��]�d	|��_Oh� r��w�~����~+�"���cx	*�M1��P��m����s�-���}�{�c�co
�vT����w�s������SN9�\u0��Ƕ)�V(
�B�
<>��=T�1�gE@���#.}���w�}w����5>�H:��Sc\.��3�Q����q�"���0$Iv@�4�E|���m��H!�gi0v0�@"I���+�e�QUF�}Bߐ4#a�P	\)��6T�1�c�%z��Nc�+�Ά�ial[|K`c��]�hݑt#$e�p"J�Y�x|q�=T�1;�v;�dc��>�1�ţ��fx ٥�h�\��s$E��|°#T�cuNA	�B�P(�VH���7�*/@�	00T����E�1��US$K8�	(~"	���t���2J�&���?�9�2PіB$rb��?$����������Y��i�NH��,;@�4��J1�ֶT&�#��^��R��ٵ���6��J�q�o$�1b�Z��C��d�<m�������l<�H�sU�N��i밃�,%�
�B�P(� ŉJ� O�d�$Fm�_lz8n����O$�1?��������Fb�3Z�|�c$�t:7�v*[�c��NFLQNՅ~�:F���f�ʍٳ��<��zJyi���x�=��W���@E�����:�zH~Y(�V�T��\x�˹Q������1R(�Q��ХbFs�X�T<sS��T~�r-��Q�Sh�G��6���m�S��Mʗ��S�,I��o��p�*�����Ў׿���e�S�IP�ة�*�f�}4ؕ�
�bܐ3kEn�R���~�h�>�ؓlI>������l6D����g��6�Iz��d�����.�(98�G����VEL�U��Z1V�Ud\}�0֎�|NM]#��ߛ�*
�tA��6%���R8�E��&F�r�񰀦�s��M�J�q,���|���u*����.��ԟ����7�Y���}���8p�����U:��@+�
z��]r�%����Ia�_z��$�[Ȋ��x��k$�>G.�V(�q��`�{]� �<I��b�)��m�=uo����D��T�DNlr��ض��RZ��
��٤i��_j�؛��o8�N�+��B����}o��9��h�X"'����j[�1�nֱ��i�B1���>DL��~K�%[)�*+E����]�MRgc�����/��ۉٗ��H+�S�y;��J�k����W]u�\��<*gDy�;�YN�;V��ԱW�k�.Ԝ�8v3n������o%�
�b: vϓ�s�#h�
l��"݋�T\�["�1��g
��S��=��J$4��Ģ6ǌ���<l�#�M�1�^���'?%�8���e�*?v�]%Њ�DӍ���S�i���J�s�����B��N���&5WRd�v�����y�X����fN�{��)�y�R�B�M��Tbi{Jm��A�\��D�S����tm��w�
�Mj~����&J�c��I.]�R^��8�Huj�B�PL�Hq�{������i�r#�Ҷ��w��Ę�9��:m�+��6��m�]<T��m�6��{.����%9Ǹͳ�B	�"
�|f��ѰԿl�2$�^�9yc��r���7�t?�y�s�՛�΄��Bl�&`;ҕ��������8���>[8���?�\�,��q�c�x�(����IK����M�S� b����'�9v��m��mR�i=%�+	DҾ��R���ұK)�M�9�g�q����J�L�����~M>S(�VD�S�}�C��.���8�� !]�m^�Hybf����3yF������mp��'�m��.υ%K��΋������I�C=����a�@�x���a�֗\��������=��sr>�b_|q�o[�jf8��~��׷8����y�,b*bS��>���}�����#Q4_��i{.p�����L=CrlRRv$���~�Yُ�M�X��u&����H��P��ם��gOֵkזs/��r�#���!ݴS�ʚ
4��H^s"���#]ƶ���s�9'�.�ݷy�f���+'�@c}_��W�Yg�՗���b�J�яA�ĉ��v=�q��[��V8餓j��v`o������z�#{1ACJC���/��K~�|��T~�F�'i;G��7�����G�~��J�K�!uLx��6�hR�c�buk:$�S��Zш��Y�ES7�&��"��n�m�.��)U$�~2;MeMű�2��W���!Pɞ;w���l�ju��S�˵3]�"��S8)�Q*OGr�1�ʯ���#���5ֆ|�~���R����)�ܦ��K��o��t4u�b�K~5�W�hDWB9��ؚ^��"WM͹�*B�\��q�D:,�D?�[ǜc5�v���hA+$�O�Jy(��I�5��9�sS���M��d/F���������R�h�/u0b��u���s�12,}o�h�X[J��s�Z1pL�C/v���~s��UBrl�̘��QFM7l�i�H�w�]ߴ�M��a܎�8Æ����E�P(v�z�n%c%Њ�Bz�<��m�5�ݗ�DK���m���xǎ���	�,	�p�R�3�����$uJS�U����%�6V��{/\x���W(�8��� �@+����ᢋ.�;�g��2�B
M���k�TT�w��-��s?��O�r�xS�)�|�������˵�۶x#��S�9�����9sF�� �����/�6��?��3�/֬Y�!��m۶r�B��A	�"
�.�ꫯ.G��$)�&	QM���o)�+�=�THȸ�i$(7�|3�X��\��l	8�p���x.]p��Th� ����`�=������+&N�͝�^������{�1��k:ςb��ᮻ�*IU<�������㎾;dK�.-�U
�B1�P��U"|U����䡫RŁDo��K:�����)��&6Z��a���dɾ�ʅ�.x>��x	*�x-Z�]�<'q�� �y��K�7�����^�'Vp���]�@��0�>���NW����x�����,�O�;cxN(
�dB	��mG��F�����,���)?.�ʥD�c��s둊�.������;Lt	�6ЇM����k���J8J0�o�Z�@֯���a ���e��B��9�dx��� �v���b���o��r1lܸY	�����.1H�z��#�tʻ��{�.����J(b��`�Q!�c��ǈ��ͦB5b�K�v&�A��%���/��G�{��?�@x��G��!ι�O�Y�f�D�Z���8F��Cr��3=��:Yê�X�i��\=���Og��/�(y�N@��u�~<��a�q��f͜���b��j{�|���������?[��i�h�7�k�{��̙3�v%ЊFtQG���� 55W�sCV�����5��d�錜��d���R�q�603̝;���)��{��-�M���٢��^>��\v��n�>ki,ɭ��00�a�_-�1/1���Ir�Z�+��F�:��k�ڱ��\�ׄex;a�6��-%ЊF�yH��E�BPbN�����=�Px��\��tNG��`8˨�i6�a`Z����j�����3�k:�����㬈��>���Mc҉S�k��gD��9���g"s�K$��.�=#��4��g��,Y��a/�ZG�m�x��Ρ6!��h�N��j�K��X�}��N?�tx��������g��o{$4W/���a����/#��׼J��.�t�˟�oy� �SU���P�����B���uʚ.%)�J�5嘄;�.��J��oR'N~C�I�����]^���L�	TZ&�m۱���B9�Z/����?Hw��r{S瀶c�� 8��8��N��ឧZ�i��'�(?�R���S�;����N%&����7�}�5�4�b�I���ז%�wLy����@~@�4P72�c)͠��ƺ�=P�?e�"��n��#<?B�XT�!�ý4�Ts�l\����UKR'lrsU�+��e�Ww�;�f�5Su�h	 ��V�m5B�K�m�ژ�=M`�"���Zo|�B K@�{�MO8+�G�SX�+f\Nv����I�AH]�?�A�"+N	��b���Q)�|��G�CA�nS�<�mR�%�o*�W���ωX�Ǝ�0|����6(7�6J]�s��`�u���S�%�� ��]�[�k�� �C }����5~&\����xՓ�������4cB�Cg<?4�� 3����%� �N�:���{"^ 1$^�Ʒy�x�T���k��mk�U{�ʑ0&�:���r��"�O�>��Ͷ	�hE#ھ��^N��� K*��l����ڝjLV*5p0��N9(��w���9`���n�α؛�a 6~"E�G�3��.j��Dy,UȐfB�q�4��kjle������0���X_���"��!���bL�!�=᪮L��	�q�٥.�����	��)�%i�0���n��F堭�cUo)hS�۩����i9���W��&������M	�"��a㎔�%)�҃;�=$�9��)aT1Y����X�#�nF�Q��y��f�`=�vX�:C���L������"̎�9Y��EN��|ʍ��>�Q!�\C@�"��MU�sbiaj��dA�mVN��6+$ۚ&:��G������U8�<P�����9HW���)|>Ww��͒��)vA�ig{.�{O��n�hE6����8ʶ���/G!��Q@۶�J�?��)p-�?�m�
+QLoԈ�ԩ,���(�_ �P!B(ٗ��"�jiA|ыi6Arp�кPgm,d��I>)�.�9q��^�X|�Wo���P�3�A�$<7$��A�)b�:sR�c����8��G��	opj<��Ϭ�*�4A�h��Q��J肦W�Rz�?5]W�j=Uh�^�uN�x�,���6�; .4�m5��O1���/�ay!r4ưv�6�ȞLeYK|��%$�0A�#�nk�b��,b�Ic����dX�	vT�H9�J�~�5Wx�%?�W#�EUvթ�j2�8V�����~�%�NB�|�6����e�=(�Vd�)Nw\��F�7�@�
���|ظ�\�o�663�?�L�����)����i�������a�YSL��o2}RL.aZ����\�K���!9MYrߙ����^�6_�p֔p�fH2`�a�M��ك8����Z*Z��}��`=���J6�WJ��Oޞ����,+�S�k7���t>��D�@	��tT~l��4u �^uK��h�1�lJe���3E`�ٱ�!�9�'�)�Yz��v~�E	�I�޹4��05k�t��sg]��{�G��H��1+�|Y�Կڗ�Z3_��p	�8E
N#f��M\EϼpM�3QL�\Tʽ���WH�dK��6�Y`�A �( �� oHJ�B�Z��v�_@��}J�����6�QxCJ��}@����(�?�v�<�D�i;Ij�d�٣�l��a:��X;��>�&a�H]R3��E�0\)4~{p��!H0nʼ���q��l�@/����(�ȾR_�=~J{^נ��=��;\9m�H�j���}��~^�������&�o7UY����؛�@�Ǜ��:&�Z���+(�V4"�J��Q {��f����$R�t_i��L)�SArr�I�
��:1LF脪�;/������s�06�R�)��~�s�ڠ\���X�	��XeO�}�t���y��pH�g`���C�X���da�9Ɨ��[W�z�V�c�+@�g�b��ow[[LY�ն�ku��O���|��~�vuu�S	��9��c��?c*4"' ���'�9�����2�H����V%�w��}�'Ā]`��D�'R��b��F��Oz��m(��}�&�/�aky��*v]�}����v��}��jW�z�>7�#�n�!��DE�97aZkƾ)��G�=�75�ٱ Z7�7�䦂:��� M�\��S�l��@	��rT�q"�9jrn8J��X�����B[H��dI�Ou�F��g��=0Zt�&��4�Y��EH�(��]?�s��f˰��"^�oQ4�E��F�KT�����i�$���b6S1�����	�^@h?�Ww��/~nb�	a�n[n�>*�1s���n��u� ��LW��G�MM��-��Iw��1��ǎ��J�}���੄�[S�E���m�A��7�9�����8�,L��d�0��RL?���x�=����A�5�Z1�q�RfM4���eIH�!~�e��G��}�rP�ލ�m2�*Gp)Y�w8j>�����F�Z�ہӠ��,�zJp	y��4?ެ, W�:�"��J����"���9y��4�|衇�K_���n�˖-��7�(�K[�l�Q�%!�0N�#�~���۷m�U���n���(`���0�<��B�^���q�<!ҵݑH\����:�w!�Z^'�.��� ���`�$nUA�s�����uw�$�Q��P]��V��.�YǨ ���O�Z10�q�iV�&�=��'�����7}��۷��͛a����d���	Hwp ��'�`]¶9χ�TX���(�3)�c�#��G��30o�<���W�{��FX��nL�$�<�j,�^l:�ϲJS\Y&Bx�<�R�2�}#d�����z���=�x�b�y]y9�VX)C��w�fb�U��1)��qSo;���h��`ƌ87Mag��)����������a�!F`'����ϴ�/�)q!r�Nu��T���1����m��~�
;�@زe�|-�Ur)�=�9�h�Tv=��ل�k�2���Ƴ�*\�g� ��dg�,���ce��=�-���P��h��_��:�SJ�}�IqU�(�w�P�b���;[�fJf�(ޱ��H!�DC���m��WU�#	)���UK:?2g�|���K��S���k�P�7Bp�z�A���7�{���
�ˀ m����!�����@�����O%Њ�����͜9��k/X�hQ뼳g��BN8F�v����n�Θ
ř�����ω}��1�y���lS(������R��_֖<��?�I����r5�����m����Yx��Y�B������	p��v���*�n�P�e�~��@�xD�%Њ`��H�����û����y���*�����aIq�y��SWI����>S0�Y��p�3��;}w_v�({(��G�˂�p�Aς;�~�/��lr�sX�Y�Ř����t,QP�y'9�:�3J���Z<��'�^�����DB]j���_�q0���_Nv��ȥ-l����8)vu�����G�zJ�QXB���lJ3cƌA�U��,��w_Q�:Bؙ/�!�9���q'��9r��<�>�n��e�]���τW��������o�ͻ�h�@_�)?'�]�yyMs�M׌kŤ���ss���2��`b���<���F���N���3���2C����J�2)���)��75���6)ߠm�[�x��S�y(�VDq�i���>���T�֭��.�.���C?m�l��o)�t����8���SN�<� \x�p�7tʏd;O;v����9蠃��{�a�l��y0wޢ��.b�[�Ϟ�{Ng?^�җ�y�7���o}���ov�Mf����{�ǲ_E����U�V�B1ع���׬��0�,V��)��Q%�d��.Q#��I&�4n���e�1�gG����i�lL1�9t��,_�3�A����Aڪ-,�6���>��o`mX󹞦��<��@+����s����?3I#Q�5k�ZJo���~KvrB3F%�t�(	��1��nMu��+��|G}4��?�c6���4�s�W�g>��,��y���ch�_���aχ��1����Ol,���n�����7�4:�8(�jB'�(�T�4� ��9[�+��Ea��������c�i�X��ʡ��S�_��X�}��zA�@�I�sEL�;	%�U�@/���dFz��:��W�\���E��R�p+(�V$!�H�}��	�{���eKD�B�GKę���
�v��1��9�1���m�S�z2�H�O����x9�sw��A����:�
�0agv���WM�6�ڵ�����,=#�%���aK�]^�W�rU�%�Pc}v/�'�t�oKH}���*���@�v�8��뗶�OЀ��Q�:*;�;��I,���~v8�@+�!=����)� �"o������&E��T~)͸?��UJ�$8�J�|�*2���OF�S"μ�}�:�c���ʕ:N
��rcK��F.�5S)� ^�t�ΞϞZ�TTF�8_�*�!|�Z&�n�1&TpMUH���)� ���%�D}���� �:���$HG�mڻg�)�&�ѫ��n	��K, Q����}������Z��؃*��N�O9�}S���9D��M�6��8"�.�E��ݦ�N�L���:����qP�_*+ձ��k<��cܯ#�x����3t#=孎؅v��
�H�����[��ΓGϛ{6%�i�rS�J;=q�1+���y{���Bm{�~��ԧL˯y���LB{SKCM�(�VD����n�ڷ�m۶�=�B
���f�&2���nR�s��?�>xq>��A�����1U����n��־�lذ}������ЗA��0��&�{ܯ#�x�G�wL\0�/�_k�j?�ݰm[����a�i83ތ
f�ę��@��P~�+�S���L���#�WX��b��[	�"˖-�����}��Q���?��6*qӾ&u�K�q����7�����ᩧ��˖-�bŊ���:�]�&8Kĥ�^Z�M%�|����q�k�+��|8k� �#��sB�fΜ�3�&N���.�a�I�xl�VذɆ"H� �fzS���Z ��}^���8� T$���~�?)hZ+cd��sw�['����(�%KʿQ�4��"K�K6�w)O
�U9�Nз���v�|+����׿����z衇`g�]w����'��X�z5\}��p���m;c�)S(�Yz�۠{PG-ED��O$S{���W�e��J#���r�k/�Ɨ�󅦙3{&,�m�DW�)�\X�rq�am�|�*�]�����i�^�J�c��4�L��Ҷ7��<S'>�d�;��(�87���_
�胲7�ۅ�/U:�>_@-��Ծ��3�к���Q�ZF��ȈJ㶐f��g�$<�C@r����!�J�c>Gڦ�is��c�w��B�P�B�d�<�E�XZ�.�|S>���ϝ���0N���/|ҊȺ�N�UT�a�یTT�C�uqǇtt*�N�m�nI�@��@+���ks�p�m���
�B�ȇө��i�RF�Ĩ�;:&glX��3�bwFR�tvt���L�v�YlB�,�Ն��lU��RlXj9�6�AT�Y�P(�� �`b+�T�zbg=�Vx��A�\±�V�;��9����rlI6y�,�O�%�*���Ę��_F4�Ov��1�ah��/؃h��gO��_��կZ�]�tiyC�Q��1 P�h�B��>0s"g/�Y�C���$nJ�:�ϙ��[1��yL8�vm7��<��nG|����C	�b�S�]y�p�M7�΋�g�<�Jh
�B�	d�[@�"�<Y3�7�1�������6��NZ�|{�/a#�����Nk�2I�4�n�X�?y�(�V�P�~��˿��;w.,X�`JC*��o޼
�B1ƠDKz�l��'��4��I)�]��)_������u!��k�ZA?!�\&ݢ�w'�h�N$�J^
�B���[���>�Y:�F������Ld�����ҭc{r斎M]���}H���qԂ��� �Yx+P)�P$��J�
�B�P(��{��Z�UX�������@��R�%r�;��4�0�?VfN�tc'�61oJAQ�~;b[�M�)�X��h�B�P(
u&:d��1΋Q���qA�X�2OC���T��ER���oHtp�~����۪������.�+A�@+
�B�P �b�ק�&$�&J�X�`��s�1���X���R��̆��ߵ����f6kF/a�������B44�ٕX{J�
�B�P(��0��(�F�f�8�� ����3kf�����9�߱5�μ+�I�n͚L�)C �t}�yv�y�(�V(
�B��cc�'>k�՗��d��m�l������`im�sc�s�e����
���y*q-*-=T��	J�
�B�P(Z TE����7J ��`"HV�fe����1t��Ι�#@E^�[
߈����94OPu����IW�P(
�B�t��G�!F�lM�r���?UN,/��4�Фyq��j:0��#�FB:�@+
�B�P�PT�'��y��B�c����h��O�f'��"�*��
3d� �8�y�%�+)�|�B�=��瞎��U�����o8s�m�^���YѭZh�iڴn�A���e�9��T��J�
�B�P(j0.¢��^���b���Y��Z�!6.�:_��>I�MKx�~�b�9n�Q��.l{����%��;om��zlH��2�4�SB=��(�V(
�B�`H`a?�rLa�H+�%�Ák	�Q�S1mB2bq��{�%�<���OkC�����o},�	d���`OK'"9�e���}�;J�
�B�P(�l6�/�]�]��A��`2'��I��p���q��u#��*�d��4�ډ�S���_��S�v*��*���m2#
�
/���,L%�
�B�P(5X�dT��ҳښ�Sbk�V�#�nse��χSS9���0�s*$#w6�.3zH�n4�j�8g�M�(V���Ն|6��kћZ��	B˃�>6�G"b���i�
�B�P(� �4A>]x����Ahlz	�ג� $8�G�7�˗K�c��9��m�3xn+���20� h���Ui��ho |�d�Z�P(
���r;Nj�S���JE6F�o�7>�[s�V���0!�䜸d)��3e��%sڼ���!� m(�@T�d��5��g�(�QC�4x3 ��S}��@	�B�P(
��-���d��`��%�����=� !��j>�	n�2�&MEׄ�t����~Ȅ��~��f���1�M���F?8�@+
�B�1c�X�x1��^0�����`��Ͱr��үg=�Y�cwc8��l�3�Cbf+�՛V�H�T�%�:�Z��6wB��Q|�ra���J�_�#lKN2vNV�U�\W(�@+
�"�]v�^���D�������_=Af6Շy��s�:��oݺup�w����A18t�Ap�'^���T�y0*I�+V��m�J=(}ȁ�	�hjC܈7�J����K�Gn�~�6Z�0�El��L%F�&��1�IV�7+�V(
EH����1�S>D�A���]�]��@/�u��+^G<��ھ��z
��L{�뮻��{�˖-+�㰀$;L�x�;��N���ۯܖ3Z���6���?��C���à�`�6�Q̙h�y�t�����7����� ��v�m��:?)d���%�
�B�HսE����-(�9�P��)��b��c��m����e(A�}Y�f��r���������p����>:�r^����>�!8��SK��cd�R�|:���hZ&��M�k�T���� ۊ 3wO�H���Ap��|�/~��`:c���dF9��I�[�|�Ú%�������cXG LÁS�P(�lDG��6M2]�X7���jT��{�K^�Gj��<����ë^���S���͒��i�Ra �:ީ2�p�̉os�[�̦M���M��n/�n̛��C�����ok����_M�u
6mF?���� ��r�@+
�"�L��t�w܉���[��1{�l8���u�{,\�PT�-�y��8����OZ�z�3W�k�@R!�s�.͔w��rn�XD�![��e��!��s?#1��Bg��D"r'��+�&�o��W��=�� ��j���w��BH��ܿ�}J	�B�P(Z��Ę��곆��s�U��ϯx�+`���/����Mq�)�z�H�����r�h~~V���l>���Sf�5N��сe�T���]�A#�e�]=�k���B_�]e2#�7�v�ךj_�|v3oT�;Q>�"�!%�
�B�h�V$&W��|*A�J��#�<�?���
�,��g�=�L�PH
qS��4�Q�E��r$D	}��%�=�Xf�5��&�X�KW��:[��_N�#
4M_p��+d�C/MaL�����U�]�K�����w�|���fJ��k�����"R�0sJ�
�B�
��~m@N[^{�S��R"����z(<��ώ�X������1�e���{,o��,�s�󮔩G�V�]M@�z�����>�WW�CIv�zb�V�L�:�~V���3�rR�Y�"������C�7B���m�I��nR�P(�V�k��Ϩ1�)=\��R�h�a�C)g4�$I����H�;�
�)#�����gw�h���5��ѥB-WOØ	" �B�#�PLyp����(���5[����zuCјg	Rg��G��j-�=a�h�B�P�F�A.��Qa��Cq�b��v��-X� fΜY��}wy��M�6u�#g��g�}\Y��.+�IJs��J�s��X�RG����V��+����(тm��OD�6�k>Glr[9��c��F�κ����mQ��Z	�B�P(Z#�2�yk� m�t����k���um��d̛7.��2ؾ}�����<|�߄իW�*{�ܹ��xM홊K��hZ�&5g4/�i6�X�5�'*��vod��S7�FAT��6{�.���y��+E�T����}$���@-���~W��'����E)ܪ�����5!�F�9x��mE��@+J�k;\mLZ�u�ڵ�f͚I�}@_�'
�ɡ��r�Je�n�S�Q�G1=�F�E9n�g:�q�uy���J��#�8�\���K/-����d�ظqc���ܶ�S˥Ϙ��&:�Ui���6K��X�o���r�����&�%���4i��k�6��0��f��G`�
>��)'�P�(��}��_-_"h�����.\|�œ���}�S�*_'қ�֭[��믇s�9F�v�x≵��	�����%g'�j.�,=�o��I����)St^;v������h2J�4�ͮ0]�o}+�7�k����s�@�������n!��S�@c��������`�7N���.=�� ����`D����Q�[���=��>I�(#[�a�*Ee��|��ez���܎�mb��j��Յojӂ�v(��*զ���n	�ʏ�����/擭�m_���ZQ���+�=��#�"�nN970^.��kG�?�yσ��>���}��W�r������_�r8������x[>��SC'�X�i������O��m����&Mi��Y�M��mK�����?�
؈�Gl�D��v�$)�����Z��&�z� ��\�:<1E���5��!�?V���fÒ2G�B9� 4�������v���_��0r(�'m+�-��z�}�ĳF��
9�O6����/�+�B��_�����r:/2��h��3D	����nX��]�&�ͿK�j9vGR'!����]H��0�NH�2���j�o����p�i�s7F����1�)v)4u*G��"�t��Rդ����g���K��dNP%�k�Kn��X[�rcĞیو�eq�5����ā	/�Z��*�EU@IٵP���[-馴<�{��_(�&
��ڵ��fA�U��Z&����U�mz� �of:�(�&%mhH�5�\]9dD-��~����2���hE��dJq�}�K����i!��)H$7G����>U��0V�&�ۤK�be�=�|��y���M��|�J$;cMd7�J������S�:|��a������s�߹�SσԵ)	2R99�c�GPN���UQ
�0�<�fMh����O�
mXB/�'�Z,�:��'�� %���f~�:"�	j��������0N��
9m;G��z[�H�Ԑk�j���3�V�֑���hEm�p�&�hmn�����E�(Q�Ԑ��*�7��8�d����6�B4=P��c$)p��)�`7u@c��T �'�l�1R,�j�Zv����z5ñ'�p��.ݳ�v~M��nK�}��c�!�����s����;%Y	��{E��@��U~���j�\�k�M�i`J�k��_�%��:�-����}φ$�eݩˮ_tO�I����M���GK�}E��AH�y·[��bh�ɽ���Z����i��/��q��Bd�#R+�����L6�N�M��=bĲ�X5�S�C�mx�Dr:Y1S��[�̀M[�[��3a�]��J��$�8���c�-�λXX���mR�i[ʖ�Թ�{���SAn&u��$�����٫Ì�;v��_SQ��Z�6]j���E|�{E��v�� ����.!� �9坤6�yXn���Lۙªَa{?�Y�Z�D��7��Т�Ǉd��;�*Jm�[^SXè!�/"����Km�ڥ�ڞϩc���T;�x��7�q�~}�vظa�>�����]�o��[�n<��0݁��4�۶m�}<��^{m�@�t�In0w
)��f[��,)��w�M�wpMo�\VA� q�.a	�}�����E�UH{���a>Te��]!߫�M�D�C�Ye���j0�� ��т�^������1��ַe�:$i?�n�����
<B	�"1r�z���K�(�k�DTj#��I�I�?Ry��؃J��C��'�ҫ瘚Յ�炖�����-g�x��G��/�NI�e延0f5\���a֬Kk�0�`2|�j� �K.�d�s��v�m�4y��o9-�=�k8�����q;���N�,n?�C+����L����4���.l¥'e3����$U�Al gpe�8�J�V�H�gK��:h�U���۴�-D��u��������A�7T��M?�J�q������J�R�q��FՂ&��{�7�Q�9b��A���И
p��:��܆d;��M=�yD�M�b>��9V�� �<��6���vf<��#��0�m����ϟ�{����[pD����RG?�Nu%1 �B�l�\G��%k̖�m�DT�0<�V?h���BH��m���������y;9)�v�������jQ��V��v��:%@��ی������ �V�	���I�P���-�A��۪}��~�!�T��m7��#�R�,M���m1�ڔ-���@:�9>+�ªU���q��׿��eL�~��W.��t��Hvr�6O�o���˗�aF�zC3g&R#F�{�|	���H�HW���|^u�������؎�CJ�4�@ʳ�K�+������h�,Wmzf�g��*p���Ƅ�
�/ۙ��7ho��a�w|���m$��6��D�z 8�����~v_+��7�xcty�Q@ۇxS�QWM'Mm�R��˔�QA*4�ԙ�V=��\J���K��L�*W^ye9+�~��8��nTV�o$�|��2�n^����أ��j��4�����湟���W��?����3`w��!�퐄Xj��L�k���,���f�o����>��Y��L�sh#�ِoU����/�-}Y���%k �M#��1 �9���<#�@ ozӛJ��h�7��&���A�j���"��Mq�MǦ�U�G=*���m��αQ�C��
vp��a�Z:j8h����5.�"DH�5�8]���fK��D�����Yh�Z6-��i���q��L�*.�yG��q��,3S&��S�Y5;*CҸ\E�\�dAW��fu�@ �jk�}���3gv���`p��F�~��Ӊ@��X�ڨ�b/���*�s���ˠ�TNl�T*�(�++������V��);�05��>È"}.j���uQg�Axq��.`�{�(��.�i�=��� �6 ��*�����e����N��u�jPw^	�@���_,�6R�q�NdcP1��Aw,��D��ц�N&ڔ��
�4�#��"�po��>F�#�1B���b�̆�h���|���,9yc��[^a|h�DT��ܧ�9�D��HpG�:@<O�U�-�@ ��99�C��V��;�{��F����A�5��2&w�хȦ�s��n��|��
EpD�*���v�Z�����~�:1��2C�����+�O��Ӹ�Y��KCrꓩ��m�g�_h����!�tR8�n�T�+��'��#����d">�����mS(����q��3"û�`�dH"��S/E|�J�J�o�A�A�l�<+S��B))�Pg��i0�X�#�x���\ZA�.�b�m����u��Ykj��u��4�	�q�7M�������EО� �����	�)�rc=���c�Su~P��m��ؚlt����V��;h�2+#�z\�%�^���E�"�*�E�ªxi�.��)B�E%�Jr^�9HQ8����u����Q}����uA��m��'�I�	�@ Ϭ\�V�	3f�� 4�a�֍0J��v����r\�EێTW"�vƇ�.���6��=��+YV(�aX��z�TUK���)����!գY-�4l�4se���|6]�9c�n�i���_�m��hD��i�f�<[�gK������؃D�aL��J���|�_`�Kg�����O�2��#�a��~�z���,�������4_.\X���{�q��;��vV��\n�K"ˣ@����C���2&+�b������ŋ��3τ���0.�����'?��N�b�b��d6<�1u�g�:�c�i��L�-��b�\VV���M�5�&h�j����f>CH�� l^�@'ĿW��lJP= �Y�
6��h�>&�X�v��L�J����y�'>ȷl�R�MpE����/H
G��v|����mǉ���.X�l٤��q��r�V\��c�;"�Pa�Q�'��Ʀ{L�i�1Y�;w.<�9�)W�,Y����D
��r�ߕ!���Z8�(M	'_�5
Wm�1Ԕ��;H�NR����u��.���UjVv�n̍����&,��(�?D� �m���oC`r�J��������U�Q ����K[,]�y�q��d�O<���ЗqBL}�!�m�"m,��sSL�T�Ӹ�\����׻͠�~ڙ�UP(���j�=��/�(P`�h�*���A�B�2��H������~��=bZ��d��Շ��NA��\mg�a>K.�C���i}La�)q�aJ����Ѫ�a������ջF�⋴b���ﶳ���)��f.��isl�2��b��'��$�X;�vV⬘09���o�r휥6ةj�|a�N����M������'Q6�jt�/泳)	��c"�Gl�V�m<�Xm#|V�;�s��p�e���@y6�F�٨P]g��ّ~w!��{?�s��؏�q!�9ǤM]b�dP�P� � �c��s6��R�S�O҇�|�<6:f�ۏCSɴ����/�Fs��㰍�G�#Կ�ۯ������O�b6�@&�Y$��_��!WU��8(6h%t�՜p�~CgƱ]��PZ)3�/�B���vU umf����R�^x�J�(jv�A7��5�գ��q@H]h�A9Igl�z�J>J�X����Z�|=��\��]��Y���{!��xv޴<�����\O�,�[���?+��m��k|�F����/���d���J�v��(��a��s��w��.q�
Ex��Z�LSQ#��:)�����OÌp��c��%�@�qFhȗ��W5 2w5�o���l�O�Zq��Ve�����T;��YzmS�mdUb�F���曰-�9w���ї�C?�*��ɂ�g�N�~^ݷ%Hكk2Hy������br�OSg����7�Q? �b�0����<��j�	��uN����F瘮
��"$��C ��3B���aG(�D��N��$ѕ�-آS����$��IpSHq��PS�]? %�Է)��,�=^�p&陬����\(b�qT��6or�v�����gŰ!�4��"���ɷ��o�+��ț.B�M�t[��	��ʜ��Poϰ�a*�.���ü��l������e��U�%�N�b�֊΃䥂���I>�	7-�[~ah�C�{L�y@�z��ʴb'D�)���E4�.�,��I����:N����&�#�.���a��v��@yF�(7/t��x����o�M-���.D��2�9o��09f��t���S{�x�p��τf��&~�S��������0!r��v �Mwdjm�	sϮ	�����e�z*��Y����.)ָ��b@YA�����}�ЕT�
��5���Q,�|\�Q1�p�+�s.`�V���*�0�<fC8R�B*;�H�,z���yC̝��t�� �Y�qdҶ	�g�>.?Qo�:_ե0qr��o	9-˹Ib/��L�d��KhNI��SA�iۄ�-�@)�,�R(�Rd'��/A"�9y��6D��6��BG-|#ן�<�F|�T�B1H�(���Z�4DS5�h�{D��7�>�}x��㗡R�3XY�bG<y�<aҎ�y��pC|+x�֚���J�?�a�e[�\���*Z�

�eSm��L9���{�|E׍���Q�K`ɼU�xS�J�	��d�S��4�Khk
і���5m��u�0L�U���WC8C�6y�-}��8�(ހ'���g�,���,X���׊	����;�xj麰�K_����R�M[�_N��{���8����:�tD�ڂE&[�֬��u%��[���C�]Ё�DN��(�$r��9$[��f����W�k�	M>t�9f#�[����^�p!��.��ޣ��75k`TV �Θ={�H�x̷m�s�΅]w�f���s=��(�䬂���3b���?<����c�D�<�0�}*e6$�DQ7!�}������7$0b�/l*S��X��8}
��R�\������|7�����J�'���\h
�t�jц��eĈ��T�jP�Sd8e_�3�nSM��7$�HP6m�4RDu���%yڰa(���xы^�v��#�� ��U�V��իa���� p�s��;��]=��~�P�����=�'�
�	�i�.4���P�]��;��iP�y������-���ӖW���?+�]*���g;�{��NBM۬L_Qf� �?{x��~�0:W�tB�+QV�H��~K������|[n�t�ה}	��,����~�zx��a˖-0*�s�=F�!�cr�'�g��<p�e��*Щ�s���ܗ����O|��#��3�<㶵�$K�7g;P�k�(�\�����D��2p��bv�b�=b�1QicSx���o>Dl?Ch��wz1ƫ�N8�/�M\�5�RA�8׊�j��fh��34����rV}%��@�(���LQ(�!r�k����A���\[m�L�@9,U�;v��7��B[_y�P�SO=>���q����K���9I�+'�|��m�7=n��^{�Dߐ�:�9�]��*^����Oi�� |�~�>����,-�9I��H�����_����AŬ�kL��Ў
c���V�`j�Qv[M�Ͱ�;���إ�M�Μ�� 	�S�6����A#���۴�/B)Z ���:���C�c��V�06��������wՇy���q'�{�w$H'�\ +V��QA�AuҾTG�:h4���()�]|�}g�	'�P�痼�%%���pl �D�����t���Io�F[�G#�����,��O�>o���`j*-��=��b%�p� v�xl�дV��H��_��*���°�;���XgP����Dxs=r<�?� DE�gR��Y(�4�>r��b���>_����ŋ�w�쥹��a�w�����fn�^z4pī&�13k���?�cJ	���lS��2����ۄ�LwR�Cx�bɳ�MD�T�:���7�qϜ<��R�s�oJ����r��ON�UtD���
�4L�db�Sp�H��J,%"MⓃ��@ʍ5��S�EɱӢ#>�Hj���D������v0j�G��tg�vĞ�_�eR����vN@	�Tbz?3wZ�9g��9sfu!��l֬�`��c� ��O�m0{VQ�0cF�2�퓍��j1(r92S�Re�*����&�����6�xg�@!�)m�$sR�ɞ��B<h�1��-�UUc[Rg��lB"	�c����i�-�)2W'!�n����]���0��7�xL��V��vX��d𞓫ADI�}lF��$w�ָ��ϵ����Zn�=Y	�B1D�.��wFR(�$$��M��d6�����VaG�7,қ�3�m6��w�}K��>��mq��ZJ�S�)[���s�R�S?o���dEޜm���<=�Zy��e�a~��w���Of#�h�1�� W���vl���
#���j6��T�È�3�E*G�5GQ9Y����v>�����a��U�$�p<��χ�N:���j���[o�k�����h�0Pҗ"�S�OG��A�hJ�%`��c�~����H�i:������c�=6��9c�%�"E���5�;��1�O˕lH!$��F����:ѵ�jә�K+A>_�!����lGc�9�f���V������X����6�%�g-��۴ۍ���+զJ����� o�8 Յ銋.�~�����(R*t��"mb]s��0�f�����}��bX���P%�C*χr����I�H��]��ca����o	��+��ڐRP�aY�j�(H|/�nQع���مM�>�#�9��H:� eX�\G�V��M�����qw9VRz�=� (��)�Ap���H=��XJUȵя]DS��Xc��aT[�>���k?��-)$���v��$иX�E��go{��-3E��X�x{�/��co%��� ��;��g��lڰm�x��F�,k�~Q}k���l��q�EX�D�]L�>'��"o?�� �g#�ٵ_�	L6��z'BnϼM\b��Ky�@�ߎ�G����&��Ҷ��su�ж��N����ʈs=��n��6
�EJ<i�5f��)4Ͱ�f�n�-X%��s���r;Q[ݠC���h����.L<}�\�K~y�k���4�g#��@���!w/<T���ږ�g#��g�||H�ܐ>�#����L�z �;o>̚0��֜3�L�<7O|�r��ML�ٔTߦ�/��R�i��S4��CG�mD�6hs�G!m[��9=��<�8����������g>����Z��7��� ����Y���T���Dz���S��b�������`�܂禖�օZ� �F�G�W�*Y��ȍ�8h��ex�����f,�
��aΟ��?�/��p>�XV�MȮ=WX₶3�Ïi/K��UY����?r��=&����X3��
�^�����_��#���!��XO_���#5&�*K���n���!ۅ˲C��nM����a����D{v}�O%��܆<�l�x�'��br����_[��̗�פH�k�MG=�,����'6p�)L���źXZ��3��]%��.�K�P��KR�j��jz6[�L��m8	%�t�8���t�t�zU~{ͺ����QT�g��ɨ)�A��ue�\�� M��; �il�*�hǦ����]H	� 0gh���o]{��$��YÍ�mz�z�����1{�ͰI�H)҃ XS���mHol�t�l�����"4�z���*J��Ee4E��ԯ��tD������ۧ?��)+������������R�=��Tl���i��'��Ƚ���$�gE�l�����SS�3��km�>��I�Z&�^pf�bJV �< �Dyu�,qvJ�	�*���>��҄��, �=b�bo�D�z����Ջ���L�w��Jj��۾/tb�b�Q=`4=P��Ɵs�H���M5v��nX9�s��rG�6�֮��J�ˌ�M�C�7Az���+�k"f9�q��.��q"�9o�(���8��8	�SO=6l(�K���}����t��)]l����yFm��D��U\˒ڢ"|V��d�F��4�F����l#m�%��Ӏ�3BRN�/Vǒr�.9��*ؽ���,�ذ}.�Y:v����ٗG�<���<�AR���]���N�qd�!�۷o���v&��R�YI�8sf�5�WɾT^즙�!�e���fڋ"u~��t��C�)�QIsҏ����Sަ^�On'��+��o���t�R8�裃��{J=��N^�Iٲyr�7�ΝƎs/�gPN	�TӪ½�a�G̲���*f�*۔4��#��t2��o�PTU1��F�r w��$��-�
�ظ���6t�v菵h�Im��=!Łφ&&���	4J8������sa��g�c�Kx��a:���TB"��5Mݤ���1-3G��%۱���hݥ;��-U��a�����s��݅4�U��ֱ��Q?�-ڒ�X�b��������?w�y'u�Q������1�:BbD8����4m뚾� ��%Ȕ�Z�h�R8+B�z����QH���iq�9N\W��'Ȇ���$��A�FX��Q'����u��Q�0����w��`U暳�3�-bCH~�Q�YX_���f{h��SNy�{�_��^�2X�z�������ye/w�"v���{�B�QJ�C���o���"��&:
�����6FY����1�9��� �t���B��u!�M��ǣ�>
K�,�W��U�|�\`A���R'���is�6bD�痞t_k��8J0	i����\* S�,�(�6���Az�6Ea�:��hW��p��P3Ru����2xG��@ר��v��j���^GA�����SH��P4N�s��o�s����'k`���g�/x���+_�<��0]p�}����i[༝k׮�a��:��6Eh�W�)խ�뾱B�PHw�T�BΫ����W������]l�t@��QA��m�J�DO�l�R�_����W�Z|�q�9Ef�s7u����X]��y�r���2^1�|9 ��6�-9��Xg��g�s_�ߢl�$���|��0v&�\ڐ�S�d|Ћ�)�VTeIa �����)�v���	����vÎF'�.�w�띥ڼu����	���ؼy̛7��wúu��������3��t�w��X�xq_7y�Bh��-�Go��z�<-ߞ����6mo�Q~�vz�K� ./��S���2�%��WB�<�Anڶ�,'�i���9��T��
_�2��=���]vz�p�G���.o3�����܇.�����?����Fc����^��X+��ȉ���i��oUd!O��r?i�>>څ~T*0�c���g��l�;	R؄d�g�R�=��`��k�Ku�b�)�0��e@���~/|�#�{�����a����jشi3�t�-�o���Κ ����K/�5k���N����oSb�ܛV��,���op)F��M�z����:qq���[��U�g²!���7"[��*�G���Je����l�:�KG�n�����X���֭[��k�-E���:>�`�1�Fڄf�B98h�TژX��K$�M�!%y�Q��ȕ�^ѕ�kD0`�l�A-v61���N8|6�O��ZRiɩm�X��C@c]̱��Kj�Q�	���H5bN�7���F+H듋�����e�USw����?>���{��������/���ϯ���;1��n��+��?>���+&]~��is�N���=��4��rU����{#���l�Q{��y��o|v�}�^�mnߦ�k�����ǆ��ܹ�m����^ ��b�
�J�=fS}��^��y8��6�>��������g�g�	�w\9��$��YR���>�j�H��( �D��E������-P�j:;g��OI4�<�1j�9�倮�V=-�x��g����'t$3`��]K�=Q���c�r��m�\�(��x�YB�j;%ѮSo捵�@4^\g�����׿��K�_�"�~�o`�]wҡ*w�?+���>����r�����N+')ڡM�f�qe���S�]N�� B@<���3��w=�_0*hK��!cm���^u�c\��0ڹmZ�����-��w��<v�a�g=��]kT��l�\�����ŬY�������yG����~.��!�D��/��R�@ȣ�v�L�sl�2ww�ܱ����[Ԉ�Un�����׉ۢ�\����BA�M���o���2�{3�������_�2���-.]�p������]S�f����>��?�ض���2X1<HjASl���d?�Υ�Sp!���k��A[Ŷ�1�}�Ϲ���˭��>Uh�a�bMۖ#}*�|^�x�p���y��v+��s9��qU8�qPz�;N�7��w��p����pBe��і���M38�lC)Xz��,�"�L���V}�|ױ��6Ja�z����>{yFA�D���0$��\ρv>xw���ɿp���E=l�z�m�	z0
������>��O~+Vԃ;�Ŷf��������[���޿�,�!���fR���j-�f쵹M�[y���Ks�7a:�ƶ�Q֎��ߪ�Z��3 ;���C�)G�Y����0J�  v�;2#��%�Y,%�<���j�����������( z_,\>7L1���{M\8E?!I�Xl�������D�7����_�_���p�Z����8��˟(c��������^:�M1o\U�l�t�~J)W�/$��b�%��s�Kh� 0���i�:*���N�V�����ɕ�'����nQF�|[T�Ծ��6B՝�2x��
u�J�Uڄ��G��c�ݢ65m�b���>��ɉ��(a 
tS�E���SO���A�s�'�-�=��5=S����(�������&۹�klnN�t??�֯_U^�}�d���F(��=}��ՈYH�Lö������iL��s�,\���`�����#�s�4��`mU?���+��l�v�
l������^�f4Q�y��kS'��
C]��9�J�H@ze-��1%8�K��-b*v��Ma��@[�oK�_��1n�4�!�R����?�b�p�rd�#�EEn��\����P��'��	v�ܢ"�q�Jwа
�h� -���h����Y�׏��S�I�	!�mC�:�˕ڀ�2lx�gˣ�!٧��P��h�j���z���P����S�+�r�/&ۇ�2��!%�u�]�aA�^���;��Yj�Ä�TB�Gkq�T��l�xeC��?�l�Ē͚�^c��	i�eLl棔��XHL��4A	�N�ԛ����4)U86�0�����u�"6�E�����Mhʠ��*��ܥc��M��
Df١�,ˠ*paUmC�9������^������$J%�@$a���&�6�����v��fq�k���ov��f؋I66�M�AH$�$��BBH��ݚ��[��:Lxo�{�if��+�L��ӧn1��lT�f��:��-�����'�W�䆪�>��l��zC�>TNP��݇P������+�o�!�Bi����w-��=w���*O-%v�B'~�[y9��.�	���=�V���e������T`LԷKtq?/��3|�G�).�VIvT�_J���|�#o�Fv!|L�F~�Be����@�!�E���0�>������p���h:���C�V����~V�� ��a1W5�>�oX�.[W�OOF�b^�<_�sc}A�茂\���4*����Dt%�1Ot��t[���PX��J���BUB�*���
t��ۭB���@�*h>e|�eޫ�{:y0���8������󋦅��ӄe�gޗi�i�3���%�i�й̭�*Y��B���(�U�&�����1r����iC
3�)���3E6�fyl�Yf���~��ܮ�;�Eǔͻ�vPZ��%�^e�I�X�Ⱦ���t6_b6���`\��G�כ��L1�0A��?E^Tj� �q���շV���d��>��1˝��ml"*m��y��d�i+!�f?O�xt ��+��������C�@�1���W���/�`X6��	��7K�ߺ�k����.�^��������-�C�~
�
�_�h�^��y��*>�z���sU��(�ͫs��O�lV?S�=�
��	�gk����!�I� �����(�	ٟ23G|��IB��^��pm���e*���Q���<V�hZ�[wE�&|�Y9��W�J+����ʨ�@yۂc ǐ���ɟw��"����݇P�k�EР7�P��m��G8Bi�:T�v�������O�M7���V�_�[o���|%<���-�ðaCᓟ96��!`��SO=�G�孪N�����߉�2��#�PWi_��^:D�;��V�LUTCh���\+���5�㔋havP�N�3Ґ?�d�*�U�!=���$_�W��uKb�t�[5�O�;�c��߷c����p��C ܯʨ�����N��ͣ��hl�*�묳�3�*uo��^�{͚5����|ƍ�?�ฺ�ҥKAFH�)3��#�E�Bci��k��S�L�Q�Fe���`͢A���:2����P�cl��p�`�͠_?�37}�
yw����2�dQ�U{��2Odb�N$��X4��"u��G�;�T�UT�(��ʻ��0�N�����n<�민gKw�yq]x�3Rkۗ�i)�T�8ۦ��#<��2m䷭$]Tż��)�;�]
�>��F�'�S����<=�m'��x$J�{���;����%�0a��|�UW���^Ziyo$χ~8s�1��Y�෿�-�k�ND�M����2��龲��,���'� ��CIt��>k��f��>�v�sb�n(;@�տaA/A�Jɤ㐔�&N��d��,�̷�*ٵ�2�F�5Kzg�b�4䓔M�X�Ӌ{o��X�L�O��z�\9NoR*U��J�����J�*��6��HF^�I���=��9ϻG-/���V�'O���aÆ�c�=w�uW)f�~���H�w�qGX�b�&Θ� �����13'�E6�Pe����\Ei:*�Jl�`�l?�$�U��X�����<h�y)c�5R��
i�I�-�?��>%�d�OD$�@UY[&�_���?I:���M�y�τn&�G�kJr�o���A���H�S�-�ֿw��}��mb�ރ���hl5��G�ݠĴP���XB�Q�+����z+L�:&M�[l�x����3��믿^x<>���G?
�o��>��?�<�r�-��틈)�1�!��b��Lz�<�ʳ��^�̳.��y�cY�A��Rw��ߡ<RtVɷ��]P�����������	GDY�H���*Ɩx��m�`$��^2�Q�I̶�?�WW�>KLIٙ[�%��A�Z&�Ё��g�l�&R��P�WrX�J�v�ZA�)a�4�;̈������8G������{���ok��|����o���X�jU�������[o�z�~����cx����@�c~Ll�a�&W���&)�|��v �-�����+��ҙ�ۤ�b����Z5���^��:�"��9�=��ݮ	A_�"����G���r��<O�H�4T�_{��,i�*����5/��l�6d�kZVH��#�ld$mf aȯ9OdPa��)�b�� hP�G�X�p!�x㍰�.����n�l�	|����O�*ɨ>�c�-��R�����|�~�m���1λ9��<��e~L�F*��z&CW�ܫm��\��_^��ֽ���h_Y�t�w�٬�e�r#Q�=z�M�{ ���*��<(?�x'f;�H��BŚn3�q�_�G^ݼ|�z(/�T�����m+��i'͋P�(��O�@Z#*���jǓ���*�C�EhT���>�0a::� ��봢�Q580j�6�l��g�A#i���;��A!e9�=�VSĔ�<E�n��:�(}�@�!{,M�Rݦ(C���Ȣ<�H����ی:�3�,�s���|M>EO$�V�����Hϖ�֕���(�13V�ap�>�׵�5���I�Q�j��J�ʮ!�v¢M�4e���l��$����l�聫����u6t�t�ɏ�7�b�䭺��l#{��F|����n���m��;�<�H=�0�#o|�3�Ѷy���_��X�l�#6a�n/�7�����_:���iz�6%�KZ�M�)�9�>����z�F�)V�f����K}"�ap�#Ōu���!�#�&��o !z��_�6�d^���-A�P3X�l�8U�F1UλI��Q�L,(�|�.��K�Lc�	�������6�z�9ڂ@#0z�=�ܣU��^��o?���+��@�F�c�W����n���z
�"�U�E���lh>��(B�R�w;*s݂�Z�ވG�Y(�67��e��eT�2�TI[�@s��XՓ�E�ř�+�w�Oi�/_,�9s��[o��������kqk����.��[�0j�z뭧#y5�l:ְw*�F:�0���[�5���!��3*�2�9����~W�%��59�#��Z��n����l�����r	�ヘ�9�c���j�)ä�@�6oSWp�H��tV	�h�:�N��p�5�\ӦM�Q5F�	'�p���������4�=�\{�-_�7������*JP�����3�G��������*js�u,�d��w��4e�ӌ�=��׈*ג2������a�����'ꧯ������ܹs���B�o��%��N�>��{o���#�BQ��w�yG�h|�}��=V���(���PZɕ��I''��E�I�} ��RK�y�=-�w���(J���[G���r�fk��ZL�x=\�k��bC�����g;����4��%$c�mhģ�>�}��C�Ş{��h�@���60������r�_��W�={6��%�n7iC�Z����R��,�/�ާz4���,=��6RnU����Ӿ�E�r=O�h�N�f��~�;�ѓ�<����f��v��H�z��@+W�lJ�m�q��O}
6�l3M�M�y����{ھ�m�=�����|��סP9�k�4�vM�j�\+@���:�7QO=�����[@�39�V_��aخ�z�S���S����y�fQ;�g�4���N�������w�O��a��PmE������1c�V���I'������+�x��O��m�}Fպ̢+�	�����������ެ�_�R�*C��l��8���ߤ˻��	pi��/x~�m0=�����vD@��E�B乑�ChwBYUi��=�j�6�
89���N��;N����'�ct*�O�=Z���6�`m����#�<�=�����G����X�"Rl^C���y/��KH`���X�P~E׏��cơ�����|��������zY���1��$��ZAL)�y���ħ�nё�� �N�7�1I"�nG��w ���1I����� x�%�7�cǁ����n���0T��;�W�ӟ�����V}�m����$v�}w��g?�u5�:�ꫯ���������S��"O�Ձ_��)�cP4������I3E��Y B�WD��U$���N�*b�\�w�$�y�{�V�qe����vF�m�`�>d�P�9����|\G���� m�z�s��V��E�>�/e�b�+s�}.�]*�ʫ�7^��}�; �1KLC���LQ��@�5J.�+��ȏ����*��"�v3���@"��d�	��rdx^?/Im��d��d���@O���{8����/��r��(���]_$0*���{�@aG��/t!=�4��x� �J]8�:W�2#���B�M����/*����}�W�p6=��iD�#XeӖ�;��Sߵv%��A��\f�Tf[���;����˿h��j����=�b/*���¼y�`�̙�կ~UO�kp�>��Ee;$���f��9
O���G�ɫ[��i�Rk�F�5���t�2�)�F����z���>��4�5�����S g��|U6�P����ye��`��ē{oh��6��0u�h;��7Z3P�Ƌ��ɓ�s��?l��_|q�.�B�e.��uS�ضر������c�b��,��j��5t]+��ԡ���,Q���1�]Y���o�*��mG�^eT�F�z#�ό�����?�Q���$����'��
5Z%�(X�f譮z��i�Jxq��mNڋ������@�Rk��e�n���F&�|<��t��=���%���q�v�j��)ildv@�+oC�=��ҁ�v�:���>��9�Z쟹����xǱBmlK��i/��"8�C�ꄨ̢}g��GL���]��cl��a�BR	x�27�"2B���e��4d��,	_u�S�n@5����H;cOA�]g^foBU/�N��/YT�Q8*�0�D��a�έL�8v�uW���,�^��^�c���2bׂ��u��02r�6���k�i�r�s�'^����{x��,(U�����י�BU�<3�&��PR"g{�m�Y��V�ٴ$V?��J��u`0�6a�8pV�e�]��~��7��9K�,���>����U�t�͢�:Pf�����Ձ�Q���z�2��o-X�j,l|�O.^VÐ�����/�����VQ�����O�2�C��n�s�kf;;��� �"�W�^���ڢQ�g���O|��o�=A��<�F�2b�w�S��"T�H3��
J��TY5���ƪ6�.}K-�A�8��y72m��;cH�Y$������㣼:�Jy�^W��!�᱑��$�n����m7��������gآ��`��J� F6����M�������b,��M�_��Ծv'�h-��O����W��3�[=����}�����!C�	��	�݉��3v����Ď�R�"r�W���9�7"���������	�w�uW�^߰o�_}��oB��f�萐S�	eBߣ�}LgژXrg7�ݠ���|��_�<*`��w�����dH$�?�����/��s�IR���3a�k��f;�jxpr�-�;W@���p���{�D�y�:L��y��HN�X��lX���0v���ů�B+Q�䇔BD��Jg��Q�c�5�G^�i9��OO��W�Z��*7�z�W!��Σungb،�Ww�s�bҤIZ�ƶ>����Z6�6ƌSj���S%����Ƿ�����E,�2���=����YY�p(ͧ\�T��3��6mHSe*6��1gӇ����i��UUm�
2�:s��di�[�2�o)��D6SG�gU6_�?ɗ���c�Z[�vJBڛ�th����c��ֶ�NDtY�v .7>���Fe��D�|�դ;��dZ~�]�bĺJޡ2h>�`��/�R��"ŹLڲ��f�-t����XZU��B�������T��
�&���/�ܭe�3�}���w�(s�T�xlͳ�ߩ%��l��J��w��2E`�T�q.K4Ӎ5��BJ�\�0K��
���|3/-�uH��$���2gճYf*!��?���+������_�[em�^�ö�4C�t	�����t�D��
4E�_,#��CfY�&#6��"��"z�	YC�y�Yt��'hO�}d�w>��2�=�⏔ː��N'�P	mFh�f���y���5:Iô���N`����D�^�ߛt|_�rb]�	h)�m��(4����j�K�{�%p��=��b�s�r&so�erbO����� b�IXth;%�^zR�&���2�6x��*᾿�_�('�Ղ�-���4�U�]�m�L���+�&�0Wy�mt��Ie:�@���&�<�B�b�.^e��o��[�X�L�J�([GA���@��|6�q�(ϼ:�Uk�<Qi�΍ ��0�E(�_�2y��s���ʵ���a�w���q`�+�M"B��<bzB��&����?���i��^cd:���b�&��(��ȴ#�Eӄ�Ĉ�f�{��!������NSKa���S�Ɉ��.��m�ɟ�`��H��W1[X�N�q�}�� �oB��uƞ?���Z�6����h�I������C�bF�����c�X���PZ�o�VA��R�,3T�X���u�Ҷ2Ş0bd|�����0~��$���W%�\3�s�0����+��3G�}#��'O�Xv�ʧ��";J�(srkTO`j&9��� ����m$_�����b�:mI18�5C6��e������}\&ۓL\��CL�ZK���&�LQ�f�%�<{%%$?��%챤"�.�n�g�ϴ����)��m�Qĩͯ��f]ԯ1�F� �F�<�ɷ�9�˷7�@���f�-"�e��Eh����-H�p��ѣG�յ	=*�I'�r�l�2�\�v�ܹ�V6*޸�!.T6nܸJbF�)b������c�3��=����!�?�xҷ�r�86�<1�}FꈟS:)�FvK���8+eH����u#�/c��$�l]�z�՟�2�Qjߡ����K�6*����׬( ��c�w���7;xI<��vh&28�'��#g]�c,��*t7_��Ū��z�B�P�υ�C��-�3Q���Ǐk$M��)��7��%�4��+�=���;�^�X���{C��������6�3��{��G��������ٳa���ӟ�L�ᱧ�E�L�y�����s���]N5� ��Mb>Z��ZK���(�)��`�H4�3[qr�g]0��˃�4���ÐSNP!%�l�U�)q����P�%v���U�'�tha%|�A��U�y�2C}.�U������Q�r��c���'FPx��~�/T7�V�s�D���9�e�V��S^H�.�G��z
��⟠�x�������(O݉�^z	�q�m��26z	=�u�"�E��� 5���U���oۜ�P�.M?{Ę�I	�%�$���2y�"K����z�|�W��>qNR��iB� ��և�(�L	�@�f���U�|X�x����O�i�L�P�Z�oS�x�{���pʨ|{�d�^�1!2�;�B�X~��ыS���cޣޢ�]Va���Ui�3�f�;�����1l+����ӧkی���@������￿V���ܲgz�X�����C�|�'e��M�R�>%�O���9�v������%a�̤?��y�vp�mp�o��LbJ!I������I�Ǵ��4S^��	i(V�^���y!��_h>Yx�M�E�L�|>כ�V�c���q�	̙3���Z=������5�q{�(��߬z4
��,�+�ԥ�����ߛH5�sp��wÖ[n�U�k����n(<�w`�$ۍD���|衇ছn��;N��̆��OJ_�����/#
�gI%�o������/*����Iڎ��8wdU���1�PU���i���l�#�AX!J�G���i;���g��)�[?f5�^g۝	�3=�^�$^Y��P�$�!�u�=S�A������e�L$�ԫ"�{\��(�n�yO\z!�KQ�W~d�簝p�5��QG��p|��_��{,XM��y�}��+�y����	���*�0a���6��A̮��U��yOCy^yOR� �n�i��zUs�'>���;F,ɦ�7�������J)��Y�@	0#���ԕ�Y�zzT'0��M´�=��Ń��?�1��JH���Φ�Z���Oib<���5�ctG��������P h���V��2*y=��)b���Y,�ؕ��h�ކGyD�}�c0u�T��7��s��wp�;<�@8����{�{ｷ)uxꩧ�7�����͘1�.���)�1{^��\��VD����z��  �IDAT����"�۸ӌ�[z��Z��b���d�!ڲ)8���"3��C�^��8��ë�+ѐ�L�٤G M��G�w���d/?�B	9D��������;_�,
	c�L�F�}�^ ��c��|d_Fi-�э)ʡ�B��#�l���o�k�g;~��_��;�	�1���b�z���s����˵o�-���w��M����x�iu@+	懫!>���Z��z�5�F�ݏ�T���#�e����W_}Uǰ�KE``F���#Y�.��K�Q��o9�\b�L���2�Y��#S���rd���*ӬD�&k�`���W{�#���P�%~�x�;{]	�i'X��i<���y���y睧�}b���_~�m�6z�.�h��Ǳx�b�5kV�>�j���͗/o�����>}��)��\H�#��d��V��Ӳ
uy?fg�輔�֛w'mw?��O��?�1�99�M��^�g�w���5���#�<��,`9O<�&���v�?^On���+V�Ж��kY�l��;L�|��l)9#��l-fB��~GsMO�Q==�E6>t���S������.��鴊d�~5<�NI&k �<i�k�%�tbD} �iΌ`B9�ÕS��S>I28�P�]�G�x��ᬳβ#K$!m�����o WF;蠃t(�aX�f��p衇)St�(�/���{�@�}<[� q?c3�v#$��g�쀢�*�M��՝���
l�_�ד�'�?
T���.�YF���12�!P�j��4x�jŒ��O���$KE������B쾧������!�!�H�eI�7�.�?�hȧ�7���`��uS	��x�{��MmʱʮɋT�;�6/O^�NF���c"��;��������dG���y] �������;���`���]�`D��W���$�e��V�����~1��IV���Ê�)K���:H����:x��ga�v�
�n��m,]�T�K8��g���h\���k�Cz1%�t�UUk
���:��C^bV�-��t����u#����m!$�㏉�_6u��t(�Y�(R7VooР�Q�~��mVW��J� ����E�>Ri큄Ƴ��:"G�+�AoC�}=� �N�=V郢�pE��Ch�:���&����_'�������zP@�	}�: *�H�q���Du=�+%�P��u}u�Fu ��'�ޜ�@��r�O�UtK�ζXo�0���ur��d��;pқ��S��2l���0J:���[�#K����*�%�:-�l�<�3���@��2d��m4];��!�U�+뛭r~���z��vVN1��g�ѭOLz����W'���	����\ a����m��i�e�f?-��J�z�C�S���18�:Rq>9�g7�6�.�����!e�3��ei��~�ĕ�uW��(Z h!�A�b�f;��f"FL��R5#���e�#��xQ��?>�'K�ZY� ֮g��ͩ�"Kn�V��2ب�̓x���GYd@-�7%Y7��Vt�3s&��=����Xa�^��@���L24����*yǈk��x#i8��@I h7�|Ɍz:�֤Q$���� �����N�>�&b@���>	�RK�2u
*㼎����<�z��&c�Žv~�"�eurq����mI�C�ʠ�'vBN}U"���!6�,��LH�z>���h�MU���Z����\�������i�{�a눺I���y�&�yi�>�C�.#�3M�X��猝�B�˦u�u�"u�@�]����:�ur�P�ih?��`���r��|�z��UPu��
�,��W���2�����8V��gs�AY"Z�Ny�t��Y ���_A57��8���l�sm���g{1$��=T捻nd���+?���gay�a��Xf�\{���_�	��<�֙����l/�D
�t��F+O���ׯ�ɹ�δcHg���B��	�M�r��W"��Z�:VQ c/�O)�y��,����C��V�Ho�L���yu.:V �*a�-�L�dK��o�Ƽ�$5J�c�$�Y����`JϹ�l�&�|�������ņp��m�xz�2�Zå�l�>Q��f9��u������;�|����J�������}���Ğo�hs�n���mAG"F|�T���y���E$��@	�Vgr�`Y�#�\%��y�ؾPY��E�X�8����E t�G9}s��58�})�6T��X&���d�o�<R9ˀ+��H	 �[��5C������ҺM��!=ۥ�*ىm;��rD�oI>��t�\?Q�֒�a�~3��kA�"��Օ44�^��f�>j(��jTQc��m���#�e�]�6�F�0p2R�y^1E��W4�)���t� Zj�p�l㙥
u��9��)�@�Y@�%�▦���I��J���=�cȌG����W8=�n#�7�u�J�TA��6u�b�r�0y��]�A ������#��=�O���}�^�,��L��W���'P��)�e�֫H��ﱈ��3�=F���!��
�#�e�-�WT�@�xd2aG��yٿ�'����k����|3���Rhب%����R�h`�izLB
 ���-	Nl��l��%����	���7m�m��/ӟ�+(s}4����S'��e<�t$��a�?���=�>|���IXg�0p�"������+\�	����z��Wݹ*.{��W�j���%����*�4V�JQ��lUQ֮!:&��g���4Z~m�!6���	�G̙J�Tk	�c���NUM�7uJl�S�!�f�)��5%�@�7|��!J��t�Ds9؞��g�N���M{ �8�d�'��z�}`7�-Ň�q���3>k�_���7`�}�^��ҟ᭷ނ��СCaڴi0y���>\J��G�ĵ�0c��l��2�cѢE���~�mhwT!s1+@Ub݉^�F�y-ӗU���9��:w�yz��JHt�t���'������"��q*�1�%b+'�
�u�)�oee*�.Ē*[V��1��`�w��{ue�*��`��
�7S���O2��8�U���w��Ç�u�y�;t��Z�I ��c�=������x�7jr�lٲn�Nv�uW�߿����_��ﾻ#�A,"G�o�I�巋��[8�4�2��y������I/�\��z��2u���Q�����cn*�XVXW�t٩n�sJ�U�1�{ FZ����b�/8�9!�-�L,i��`�ĩ�佧��]]���/i�l�PBm�H�!�G�T%�{�v:��s��Hh�|`�=Z<�=�N�)R�РA���G�3�{z@���OQ�4jϨ�'�	��$T�V��U��ޗI/:ԇ��%a��y�r��P�T��hG%��x8�M�&�N,��tՑcS��i9n�eҎ��wNF���,I�� ��\Qۊ�����3��Z��$^���?m���(g�H�6v�G�S��CP?�D��S���<r�ɏ��F���ߨ�R�{��v�}���c�h��C ���o�@����K+Q��%�g]+ϑ@no��f�گ�~��u��J7Q�m~D�������ڄ$$�k�`�WT���N��%�t���x}�:ԉ�^�!��Z4����6����^!ЂnA�H�U�6RN�����(�h�����]缪]v�b�H�@ �}Ө�A�l#��礖��]����"S͏օp;F��b#�Ղ����.NsU�:Qp�q��J��Τ.4�(�EWHq������� ī�K�υ���\�����9t�@7y�ZoC�ژ�PF��+Fy����w���{�`�:�Iw��{�7�x#�#G�j"��kժU�t�R4˗/���Q�`����6� j��*�w�{o������!C�äm�è�&f�����s����YP�_�(B���j�)YFe1������ڽ����$*�rj�ϊ9�5$���������.CQ=u����
�d���ی��L$�~O��M "<B�v�c\��@t���3�<�'6�y��u݀އހ�����	J4ƛo�YOr���d�tp��w���t���ޫ��
���*tw�1c��AS�L�w�V��� k�w,o��p��`�ԭa҇����	ί���hA�@qԉ�.M� `�2� �PeHg,OQ췖�N�l)�r2��҉�b����L>��"���ĩ����!U�C�%�4[�9�L�I����+��4֕,��=��Gݝ�}Y�x��k,Y�D��P��N�]���ƹ'<O��u����9�0���k�d��X>Ƌ8p Z�Ǝ묳N�L���t|��OHpM�fa�M6���@���%4��D&�9}�.��W	K�-4���\?�2�H�*�^��D�H��FX���,�z�
�a{�ji�MH�f��#h��DY��r���=��A`Lb��#��DU��z�`L �$=���oՌ��c�-���#Gz��Fqp����K������{��;�*�D��0����5��������&	�彷�ҳK���^9�d�,|+'ϱ9u��	9�W�UچP�c�d}�.|��m�Ra�)~�D�*�	�380!����
����d!a���r��,�,:��zD��D��!ݽ����5i�0s
�z��o�c�=��r<���-!�;�#�p�	��{¸q�J)�|�J޽�Ȓ�����ܹs��-�e��8�#�⊻���6M�deh��Ld��4�]���U�/�FxD��NU[0���3����I�֚�%����멻^ՒL�v��� �����O�t�BWCN/�H׊�G��(� �BhASQv�_h�!��@ �馛���o$w$Ҹ��'?�I��k��+�����7�|����_�}��':���a>�ŐB����<"N�3��SU�ʄ�2OE���A��WJ��>qe��|��UȽ��^Y�x��Ķ�eM���G+�g���+��p�t�ʟ���h�<��!f�qy�~U�Y��XL�M<Ђ(�VG��9�\��#$[ h��[,�.�O��w��Q}H�^{m	e���Ӿ_�yl���z���/��r�eb�Gy$��~��Zk�:&��Va��PzJ�9A-��i�XdvQ�iz�c!��r����8"����s��*sϵ�%�>��p���X���p�����2���@=��N�eJa�?X�`�)��!��L�^�@ (D��X���^��љ���/�m8�I�V[meI��ѣ��c�ՑH.����&0c�hAe��{J�����bQ��:�H���A�Ȇ�{�a�^��ϴ~�KuQ�'y�U^�כ�bB6zk�Y�;����V��Һ��mQ�C�Pg3�=��>��A�Ω2�B�	�G� �p��*�J�@�6����n#���z�@��f��r����#�8��oh�2�觞zJ�Ѭ�O�:2c��pм��[�T�|�U8�u��'��hF�f���U~ysU�1�o��UUn0��
��ؾ�g<�\�*��놂܈"d�C�=\Y�6��4�Ue҆�:DG)����QO�-�'h� !X ���G�h�������r
L�8��M�_{��4i��nֺ��e��,y�>ت$=V^��a�~�<�b8ϰ2�'��se8�3Ct�U��Cm�9q9��ǔ�ߟb䓫��J����vިL!�����j�3ډ%`z�"�?RU!Ђ� 6���	^y?�*������|���mW_}5��p衇¾���]w]]C�m��f�SM�'|���Ig1�ʷ��-�S��z�U-)5.�b4�Z���1D���l��s�� �B	�V��4_�������Ϫ�t���3H��%�r��G۞S'��l�hA��]��Ѕ0�6�Z�L�@���F�4�~��'������#?�u���z���w�]��C�Z�bE�|p""h'��}18�O�,�ʊE����ݗx>�{Xf  �ה�l�P�Ԋ�OIv C��+�l&���U+y;�)K��U����+�dT[y0ۮPsy=?��N�[�O�F��i�\���CPE�ж���|�c=�	���%'�*�����9 1�yV�*fΜ�'�b'[o����Q5�F�@�s%6GU��p�>�y6�y:�ؽ V?��R��׸U���85S)G�)���i�!��W�I��]I���-t�T��u1��fH��y�]�к�yJ�9)M��E�Y�_�Q�Ccd��H<G����1@e�S��:N���l��$
����#��ʊ��8*ݹ,3�&Ǚ�n�`���ݏ��֢�4]�B�k@��	&h2\�@��c>�,!�JIp�[B����U¤:D�cO>�
y��Q2�PB�ZvLX$���V�u{,�&�\K��Z�8mjѠ��&�����	m���U����:ZWsL�>�ϖc�NJLeI��\�����L}^=� Ĵ/a�l�
?����X8s�o�<���}���:̚5�.����� w�qGf�X�k�@��(CN� N��lc�Eu�E��K����nȐ!�����5J#ʈ����!/�P9y�t,���3F��S�W9���JS}��ԔK[���?%Ծ�����6?C:3u4G2���˴\�b�[�*�*�n�N�]�LOdv8Ҟ(�O���1���dAH��o�O\?��y}�z3=�ۈ������I��@,p�X����'�|R�	��C�p�����<��b�������U�2�ns`�<��1f�0�!�6���"\D��y���\�>6�yO_�v�&�F��L�bY~�8�|\R���TG�u��y�Ҵ������2y�!��>�D����l����$WO�Z[?>��Y�ީ�ry�.KB��@P�䵬=#���5�O�no��ʕ+��Ud�Ԯ�/_K�,��k�dĔ␪ˇ"�K͏-�&���B{*�}%*�W�ٚX�k�("'ӯt��k6'3��ʵ�%�)�����	�z��U�"�r�Z��R5�X2(1��v���K 9	a���uSoQBf�quJUlc�`��#��7��M������#��@�$f{_k7�5@o�o/�˗��C��M���@���W��XT�q��E=sD�~�mo)�"\VE�y���С�B����#�1�����$��!�E+��X"IH��\��-9TD�U�+��Q�����%����>��ި9u�Y2��i�M��Z:bJ�F	'�-��֤,ŶX(jiv��$J���TL�=�Fn�b��2�P ��9���aΜ9P���J�o{`%,_��:��Wᙗ���C��K/�}��,��sD�DW��/�����$D���[F=.��:�G�C��ʏ�Mmy��v�܌L��ҩ7�Β�Yㄌ�a��t��M�{\]YZM(-	u�٫'�#�_�I����~��,q5J����78�:�3��S�ir3h����l�"OB�֏ x�cO�D�A.�@_v�e=\����SW� �Q�F��#����^^�hU�ٳg��O?S�Nu���s��S�C��P��41�t�wq��*��k�Kx�lZo�r�[�+%q�;��(�iB��?гp��[eZ�G��{[	�G�Q�k��:�z�T*վU���������)�4S%�>@0�@{.��sv�o$�Ch�@ :�n�)�7N�k1����QH���n���СC�i�"r��e����Eިb��T���r�;2��YU�[/�+O�Ҁ��*š:��mg��M-$��y'�A
���"�'Vg���Oh�POq�n�?d�@ 
�0��6�h��8�}�Y+�����o׫��������y���
	qy6�p���V�)6�g�	d�ͪ�Dz�
��ӻ��#���˨��g��b�����\���d�h!��@ t(6�dMxqA�_���9��1����a�ر��V[������{���w�4yv�"�&�A�{�ի�� �N`�*�!ۄo���`���m�͘�����Z�r�')[�j�wd�osక#��lW���ee��ZB��@ �@���p������5�C�'6�}�M7�I�_��aҤI�E�(�v�}�|B����Ģ����Xh=�_����`uW��d̘E�D��&�1�2C�!K�!��ݬ\��/t��1>֯eҖ�F�*���Uk�v7v���a3F�<)�ޞ���#϶A!��@ �0��|�a��q��Ǐ�+�b��f�ҊV�k��VOH��'>3f����B�q)�1N��<S�	�5�b6�1y�Dy
�9)��
)�����Rk%�U�D�������=��xZ�ol`R��F=I�_b������|���Lb'�H,$C��"�* N�L"���$ WD�����d���>��hl��&����?�0�Y��)e#����[�g��+��B��u�Y��EZZ�������@#�%�~����=�Ig�>���;ou����_{�V�<E8��y$�쏡��<TG��x� �%̝Hh?$l��?g�w�d�k b���̀$`��7�?��O�3.�2d�m�3f�~�h�"��Kt:��`�@/�ܹs�ߠA��Z"����s0�5���{����Üx&�Bȥ���Y�f�sB�ꔽy�b{ �4Gɡ!�[��y�|�<��Hta>&-���g��e�KFf��ؽt?�4�.!�;�m	4��4z�h��(�"����R�@ :�>�At��'^p�p�u�i%����h#�[��>�f�^K���]�H�$��12!��>�!LB5M*�]�CtQ�EJr���f����l���ɲ�{��{����O#md��(믿>����Տ��C=?���t|L�@ ����%�B'��3g�}����{�^~{ٲ��.�A<���]ڛ���4?� �X*�X=�N��7�,1��!�7�j�T�ߛ�i��ښR��,�ږ@�"σ�-9b#"D�S�ϟ�?	�@������?���mFu�?T�W�X��>��#��r %a��4���Aų(R�i����hch�bYD��� ��29S���Aߗ�IؑQ8�ΰ��S�*��硹�~C�f�&�Yρ��*�7q��A��IF���v�$:�#��lX�g/v=<��\�o�K̓lһ}t]�,1v[0�t��� L��V�F��裏���W:O��C�`�Ĝ9s2���@ �PnZ>q&�J���������*�B�XbO<Wh��Xu��M���>��-�g��3m���\�s�"^^�r q���a=�ݶMa\�*�N�i��`�w��G@�>�����^��l;6�,il;>�:qCa }���sѬ�H�@ t��U9���2-�Rs�WS����[RM#qP]4�/49�h�`hq�PL�G:v|^�B�y�m���0X��H������\���=���ۓ44S������@��px�1���{�?�����_�Z/M�۱�·��-8��ca��:.�w��]ڨ��i$ͻ�+����m��V��k������M&`
��O�>�ސ�L(5iH:{�=ΐ옪J�ir'Ǳm��ry�i~<��y�����L�W0}�Lz��4jrڿ�l�����`����n�˅�gkQ��o�kR1bq���|FH�9�蕙�B��W^y���*M|w�e#���Y���G)� #	?���a�����	��_.�Y }���"(��ZRI�3!\���t d|���@H�jn�(*�h�.��\�n��rc��mw���%�z�|�f
8U��L�
�!�5�w�P�Ѻ��~�i�WJ�@�*���K�gk�+Fm���zըiӦ�*��)��СCubz�RaLQ$�8 ����[,��4�0�� ������S����x�zg��ɱ��m��B����L�<�F�{����f���5�Z]�Z����q	.��G��v[�����CGF�@�}�'�pl��zU���[I��ٗ�m����a�m��0��|�QG��?�^{�X����L�2����镭0��7���A�A_�^�2:x84�����v$���X�= &�9Q�|��G�~�-~��y���1�H�|����*U�3�38r�l1i��>�Vh֋�Ɂ";m��y�mQdR(�~$`�xt���q�Qy�c�=���瞃/�P��",X W^y%L�4I�	.������yM�1?z�O>�d; �����a� A_��`P;�!�v� dJB�|z��3b�*O�I`�� vD�.ؿ_�]�l��~��!�g�:}�$IaY�rrcD��iLQ���c��v�s��b�$�n�~ir�=�F�AG[8F��-�r�n8F�����m}9j�<�I4.�o�ԩ��}N���r��Rc�t�A��0��1z�@ }���a,I�"�Ƀ��i�i5iȤ8k)�z]���U��5G'��_�C�U��)y�c���:�z�iiv�r�I�#j@&���<�e�v�g�-a��)u,�F����'�6/^W_}��{��w�/Ufc�@��`�������t���Q}F+�ҥK�/�����?�@ h[(�#˕\�R)B��*�xj&Um�c�n+�J��/㑦e�E�:�<��EJ�Ig�[�S:���D�i<U�bʲ��Z5��D;EGh${����+_���0����.���
'�����ZIF+��C+Ǘ��ex�gtX?T��_}8��Su�$����?����@�@ �*�Y߯���R�-9>4)��~��(�gۣ���9�y�����>����3}G^,��,��h�k������Ot4��i�MG��8��d�M��O�$'�!!D���O?�<��m�o���/|���HG'��{�&���̓�����ٳg�@ �$�rfH48�%]	Q5�yg}���A�	k��Ҵ|[��P[�(�!����s����f�%� �_iy$������(�ğn��	�l��έ���a�pR܁�?�g��K.�;�Cl�Mc�v�V��#G�g?�Y����aɒ%�@���H�o��v�@������F�H|��f��Z�$J�ޜ$>I���/�?�ʭb!劬���m/��]�ܙ��O(ѥ�-�N�v[��2E=���gDG)Ѓ�O��:��~^�h�^i�=_��*ͨ��+3f̀�Ç�7��m	5��|��p饗�^�P �ގ ٣��j��fZFT�> >[�a��fE��d֤��(��+���]�
hj�����U&CpI��~�?�	��k���Ϡc46f��vӱ�G������q�E�e�q�-㷿���qL�0&O������r�<:�@ }y�aTg�=�w!n��V��q�c^q�V�p�zT�*=��W�#[�!#�&p����W6;<C��KT��1�	C��g��1q�1V�i���c����g�}6���K (Z\0z�Q��/��8i���@A���2Jm�d`�Ţ�/7�^�F�\z3x�� c��r7	�h��(~ )�� :��v��O?v�}w���H��>�� ($��=��|�{T��@ 0$�	�F��I�	Q��H�����y�=�I��k�5�I�Q��1�o#�QO��%?U�)��s��+յ�Y1��cX�ڂ���K_��^���FO/�n���z�0p��>��N1#\�σ>X[ap��@ �<��F��NZ��I�tœ����>Z��(�]�Α$��E���p��0�������vC�wq��V��κ��vd,9)�V�}����}��I'��m�����֓��-(�>�u�f�r#YF4��X���O��C��� ������"|�F��A�7��G��k���C���l�\�ϡ�yy�2��H'��Y�_��L�}�{=7��+ mM����u���E��g�	o��6�aȐ!z��v�I/@�$�g?�������N��;^P�;�����@�W�|���W��aFDME�҅0�?��[�N���������T�g�>�`�&i�dN�� 5��h*U�,mK�ѯ�~�r��0$�H�^~�e�����k���^0��?�9<����+����>Z/��ip%�?�� A_zrW'�x�Z���#�G�C<�(��$�tK��'�7,yfd��g���mrۉ�9Q.��E����3��%�h��%�1�3�k��F�wq"a=�%�/^}	�:#A��αqi���o6f�O~�ݟ'N������q�3g�@ }I�=�����I����&��p���&�H|g�:Q^iސ�eq&���o�#ⶋ�AU?W�2��i��l�� نl?f>��M���׶If�\<��#��;��}�sz�\_Y�I�������h���s΁7�|ӦY�`|���Ջ�`\l���'���OC�Ik�^@?�D�X�`�P��3������"�Pj4Aޤ��f�l�FeI��Ǣae��c�n��e�����s�J@��v���:La��qZD����r��F��I[ªU+a��~0u�p��_��{�~�X�l�����IFF�o����4�5�Cu���m@_�q����7�py�g���?�-8����������G?���>��6�@ (��0D��YY��:�ɫ�eО�"k�X�&�\degw\��x�� ��ɷ��6ϐ"M&�}��M�'9��r�kʼ�6G��=���J���b��O~���/}�M۽�8ԕ��̘�W�ߞ��/��
���]	�^z̜��X�+����^�I]3����!�������,�;VP�?�|��{�Ku� cj�*��o��^�樣���<>� �A_D�yT���lM����n���o�s�{ˇ�䑙k!�f�=^�2y��x9&I��6{|N��x���T� ���gLy��X�M#Шt~�C;¿����>{�;Ѧ���+�t�M��S�	�~����]v���I����~�=�������D�Z]�c{x�=Y��7ވ�����?���Yg�n��t䎹s��A �i�D��`����Θ�h-�ŝBq[�,Yb�a����J#ez�)��Ў$5P��乌��� �@�͇dh#PX�sB<���8h=X�^9	Ig�i*�Gi�,��>hEM�\;��]��O�~WO������͹���[l\�������o
�ƛ�A����� ��k`��w��'�.�Z���S�h���p���7�dc8��u��կa֬���b�
�'($�H���w_}�q@r��j�F�����p�%��x�h��k���o��z�B2f�x뭷���A#��㡇�'s̚5Kǆ� 6���'a�w��/
�7���_A� ]%1l5E��*����e���Ǭ��'�~9���dg���I�z� ��I�e�hKh2�Wm�Qn�2t��K�=Ֆ�{d��̴�>2*1�#�|F��X9k�ȴѕ��a�C�c�����_�R{�k!��̙�ছn�;��̙��$�#?�J��ƍ��/|��������{�:Px3����ӟ�4�1B��qr`̺��v\�#wL�:�[o=�J�O>�}�U>�1��~_{���^Y1R����)$���=z��hP�X'�	^��"���fY�A�A

V�u����L�r:�g�%_���#�&>�/a�[уYu�{�E
�_�n��a�D��T���"� ���B�	N��,!��Px�o��	���h����|_{g���_~�����>����v�����N\�#E��]$z�&ѳg��|,]��cܸqڶ��\p��]{���_|���K� $�88BB��C�P�S�-���O�&O�N9��-�6�!���}!K��yՄ��)ϵԉ�7dW&t�2Y��p�*݆4;��2��j��Sl�s��������Y��k��k��Q�C������iUb���f����S�y��oR�9'v�CE�2�0�~("Ш�K_�����E��w��𳟝���E>@\墋.�y������sZW~C��?m'x����KX8��ꫯ�������k����� A�~�����B6��Ty�fMҕ������?����?�	|�ۧ��?"OMA�-�>�Or�p��o��Rk��x�[B�RyIB�Y5�ZD�'���X"�l"aϲ�iI/���(�v�x�	ͦ�U�:I�jG��R���m���?�0y�3��KG�k�*����/���v�m��y��Yg��#>⋏^1Ą	t�Ң��+����	�;v4����o����g�}�.]
�r�I3�8���h�hh���/�:��t���~�_�G?:�	E3HlA��7iep(�nX����c�F�5�g���}a��"K��l'��)���a�ta`�8��g\p����S�Ȥm�Q�l{��D���|ږD�ɹm�!���Z5��\�i���s�z��k3�?o���G?���B��A�����@g<` L�>]O��u�]��2TI�Zp�7���ު'� ���[`�ݧj��ȑ#t6q'�s���.��"=8:����[��&���?��{�f���"��� Gc��<Z�=�� �&����4DSU�2�)3$��	gd�_�Jm-�4��;��k��&mI?�g)	W�n	/��hM}��#���*C����d
��e�6�@�YY��_�mlg��;u��a�%0dި���j��uh,|ʔ):�V��/�Ke�]v�E�H�Ko�v�|3m�45j����Z$[��r+��~]z
|�CS�D8Ag����_M�=����N�_��W��/�@P/B��粄6F��X�$Z 4�ѣօ��'�=|���c'=/ːڬ�>��=�����D�*p4���D)?�U�yM���9 0?u�e�'��k�* ��M��~��x��qdw�͕�q�F�~s��̙l�5ٺq��V�Ͷ�	�l�ȹ��7x� ��@�$��c�t���2N4�P}>�S4Q���:0d�H{ꩧ��;����x�	m�H�)zj�(��&�ʣ�~�_zi.���"8��O阽��?�-�E��
�AA�'O�@P��;�+������X�O�����3Y3�������q��9��>�\�̄9�TRe�'�DQW>���]M�v\䚘�4����>��Tj1y����o����ķ�P��7x��+�D ��uh�@�D��oi%�.�}���*AqRUg�-��ɓ'[�1��,Y�-8!�N�w�yWt/ �o|���B�9�(��7�9�}�Yʢ�-#FzCv�"���:���`�0d��tK�6R!��j+���0k$�\��J�)��֟2AZiRg�M�2:G��-�Z3���X���zya�&��3�xМ��m��-\�ͫ)/[g{}NY�V��90��Kc�P�>��S�ld@`�e��b+k+֍uh�h�Ι\���A��Z����h�3�M<L��e��6��;�Ѝ�����eGtY�(_^σ�U^~U�.BՋG�v�}k`��ׇO�P��A��
�~ϱcB����~i�@�:8U���p:Ȭܗ��TR͵\QM�p�����y��R��_ G"C���^�r,�#|���c[W#��6Q&������ �~%bOEVd����X%�V��h}�k��&>��U�;�fC�;&?Eә�w%E�ſ�ƛڶ1f��_(k\|㠃�7@\&z���v�6puB���{����Xн�8l��ö�n���Y7�t�S(TEY[Fԣ�XA�0d�'Q��:��q"n�\RXr����*��@��Ćԑ��*��SH��ǹz'��K��,-m+'ɦA���|j��\��E����W��g�w��M߯�UTp��[.X߃b���sb�&W^?s�����M���\��*�~��и�Ƌ/��	umE���-��R�qz���:f1��pA����ۂw�y��u:Age���_�ʉ��k�ꉣ�^z̙#hAk�g�(R�A��"�W�^O�<�a=Hg�V���q�X2!Ͼ����-�.~��J�s#�3�4�\��m�p�hc���uB���\}�<���0pi�g'���?�pU�yZo3��C>�c�:����@#qD���!}뭷�q��E|��QG���@c���_��׺�3f���W�l���ÕW^	��m�b�{��>���u�����"�jO��s1t�P�ԧ>	�{4�Z�
~��_�UW]��
݁"��Lk�@ h�3kB�!�c� ���\��R�@yl�_	#��4L�4o�*M;�S�ʥ$�0`�> ��vB����d���jё:&�(�y�m6����[�o-:!� Й���:8
�a�~��C�����SO=����&�t�����|~���4YB��m��3g�Ա�Q���-�+��
w{�p�~����E<0O�@(�\ y>��c���}.���x�2(�� ��Y �~8^��m�7�f�����eH	8ɚ��(i2�s( ��:�Y�D K���*߶@BdX�N,�<���P~�V����g�������a��>��{�|�&�Λ�n#�-�Uv�����d}��93�L"�H��9�\�c�=�
�?���`��p�����H���1|�C;�W���q�)�W}��ӫ�2ޝ���|?�0�7�e8���i����+@ ��V��"��M8��En#��f�� a~f��e��W������^�H��c�7 .�/w'��kHidm<�� '�B�<G�y���D�H��&�A�|y*�Eʋ4�rk�$�d��;��~�0"Ј�3�����]D�,�p����,�����c�"��C��J����?���Ӵ���·����S��\ ���[[r��~���O�矟��]ʠld�*1�A{�*��sBT�,�T�q�<9��֌ ������4�t��iYEW�Z�0�ʺ"�]J��z�9�f���.�E�-V�7$6V~�����>=��e,.O��e�S^�6L�W�^��*|�߂_�����F�g�H�9PM����W^��Q��:u*q�a����j{��pź����tZ��ܹ�s7a¦��~�i��������$�eBb
��BIl�n�i�qX���r�1�<,UT�e�2��}�LM���"!�^r+M�ي�g�^�6�>i#���;����?�� (d
vy�Ϧ�]�9u��Q�\��/L�Ђ������\s-̚5�=��m�]a��=`�w�+V�ER/^��q��]K�G���W_���:[/�`�B![\���Î�Dq�v���Q�&��W�@�:P��2O�hR�o�'�#�ҕ���}�D7-�s	���X�N�	Տ��^����{[�/S�Z��s��:��cd7y-QN{1G-�S�U�Wg(8G�ζ�bPeAM!�|D���O��{k�'����2N����0�H�v��Ͽ�y��d:xn����91�3�F�P�f%V��	� �c�U#�d��Iba�8%�aÌ,�|��83��䗩Q[�CZ�-T�Xz߯�z�C�R�:�w���:�p�=��������}��6�Ė�V*��:+Vg�yu.H�R4	�3E����.��
��?���D㪂#F��o0/��2<��S��c��ҥ�A �'+��W��s�9'��)���;�����O�'��!�Ki�r鱨���cNt����4���fs�QQ�Ҕjˣʭ�L�z>��iq�Ӓ̓xC����U�XX�I=�}�Q�t���z����	[o�?��@γ�`��>`��mje��'�]�yϜ3�_�p�W9d- Ю�Ia�@ ($���h���
��sZBlHR�p:o��gXbG��b��0'�N�E`qeh�h֎�yy�4��Ѷx�$��m���r�K�?�6QRKC�%׶<�#�@�s����Q��n�����!�$��E ��hB�髗&c-qQX7ә��$����@�@ �]��=.W�=�x�U����3�nJ~�'��	�~�|E	\J������"*�{������n�:N&0[�UL�
���{��(�n�a��(�~�S?���R�u1�$Ύ�Aɳ�سQ�8�﵋�_Zg[3��$0�9-Է�t��X�h�@ =�Y��倒� ���q�f�O��3�l �(xy��x�!�	�"�Pu44�ΑAW����:��6}B�2��G�Y|RN��o#���rm�촟�c���>�|M�6�{��񦮴/�` 3򎳉�6�w��� Z A��Z	���2@I�w\�:2�hӧ��
�<61���ttb�!m�I�[>b���w���`�"���,*�iF(�<��gU�/T7J�=P��w}%��=����R�V�Ύpܘ*���R��Y�Ĥ�j,Z Ab�����⥰��a�2d����ׯ_J���(�GMLY����}����g�L~D!��|��`�5������,�Dj�u��=?/��ɳ#��;�rZo���և��x�Z½�FvB�i\�6�H����-Z A��7�E�^뮳6���|S�a�-a�� P�_����-�����o��Ͼ��o�1l�͖0D��a�W���W��B��@ R�y�e�'�A�@ �@PB��@ �
-�@ T�h�@ �^˷�f���[o}��>̚5^z饺�-�@��1`� �1c�|������[o���/Z �@.2v�X�n����$	��h���+���_e���1e�X�`�=���
��@ �c�+���7�G=(K�i�>7�~B��@ � !�� �eI{+�PB��@ �`�k�	lR�S�!Z ����Թs��?����v�a:��d����+�u�w�}aԨQ���:bԌ�{N���c�i����aذa�˼�V[�.��ӦM�����̈́h�@ �>n�x衇�_�j�|=�P4h�~?���y`=n��&�@sU��>��~���=��+V���V�^m�1��n�A�e���p�G�	'� �ƍ��Z!��@ }HH�y睆�X�fM�<��"���w߅�/�~�ӟ¢E�tH�q��U�4�^�t)�y������70}�t��-�@Ї�,k���h^ƾ��{��\ ��vZ.��-�ﾻ%�Ͷs��@ �Ch�4��bk�B֎���%���\��̈́h�@ �>��>&N��ߣ����V���_����y8p�����W��@��#,a<xp��.\�~��k[�:t(���:���j�3�u����5tm�ɣ-�@�G�#T|����:����>���qh����C��I�&i��r�J��K��
O?�t8��5qY*p.����f��߿?l��Fp�!���G�'O���7���9��GyDi�JS{H� Z �����zV#��ǉ��]vYf;�E���SO�c�9�F�@`;$�{ｷ&��_~9���k��i�̀h�@ �>��J�9ynt<��{�_|1�o�ȑ:�4e��в�+��C�{̘1p��F�o��C �@��Y"ʪ�!ҍ��_}&-nG��wF�G^��>��u:����^L>ʹq��@ �c��zA��y��U�70��p�j�;&�e����N:�˗�Uh�@ Ae43&r#��z��y��ٙ4����I�e����~Q��@ ��,��"W9�*ø8�&ȁa�6�|s{\��X�!�,
t7a@k�5 �6��?�z?l� <��������r�X�:�����+W�{�w��XK�[��} �,_���@ ��!��P�C�1�sHF?�q�2��:5{B!�H�ǌ���3Fu}5| �:�F��􇡃�w���@��qH�q�|E���@/��C�d�} o-]	�~���/z�X�>| �Z A���H�f`ɒ%��M}�y�ȳe����y��y�������qCaܺ�`Lq��#���!`@���7�����+G��$ݯwҮ^���]dz�;t���7����]Dz����Ů�Y�.�����@�D4B�i�f+��e���<��I�"���#�vֆ)ׁ�]�yܺ��ߨ�����j��&]��R��TRۮ�$�Q��֟���J�Ҵ��kG���� #���]�w��cѻ+�.2�`��0g�2xf�;��K`���@ A�Qo�f+��.$����$w^lk�DX'��<e����Q��F�a���]C��;6��5b�7:⛾���J������(j$�H�������AU�����`�������E+4���ٷ�9K��Z ��^4��
ϫ1bDp�|���P
"/�s��(�%��ص`�F�n[��	�����C�������@�p̫A��$5��=7����?2y�d�����F������0澾�~�-�멷��7�3U�@ �ʹq`��P^��̛7��zk�����^I������p8p��`�I#a�.=r�i�����u�2�r�1vX��7�?{o$�q�~���k���Oΐ�cDQ�x��Hˢ)Q�dQ�%���eol��7����v8�n<��]���S�ײ�-Y4mɺl�ERś3C�}�LO�G�Qwa�'�@"+���������T�Hd&�_���f�#$]���e���	A��;��v�jǍ{����Cx�����1�����"D�!B�z�,�+r�f�944Ķ�s�d2x뭷������,k��uE�� _����1Ĥ[7��E�q�[y�[�̡����8k�2ñ�ۢv�s^���[q�amRo�խ�8�"����om�}7n�oO�_^��K�!B�"D���x9X��_3H)� x�7V���i�����g?�|B�i�9ȧ4m����oo��셏�@���c�l�7��E���8b��[@�,�àMr�k��ر0��6��$���
>2��j+���P�N�JkQ�!q�� vlO`�@+�~�|m���+��"B�"D�A�]�\)7v��n�O>���X�Tb觞z
�<�+*B|��%|�s�Ç?�a|��e~�W�'�=�I�̭����[�k��mpS<\W�dy7߻i�#�ք�t�m�օ�t�:i!c�4h�&;Y���{oڌ���2���۴%B�"D�A��/�����߫J�ٳg�/}	7�p��+!A�������������|�*\3�h	4m^rӞ.�������a���b��["QM�5�Tãr��Y<��Oڒ���5kB6zKW(:_)��M���Ǯ�}���w���3�s:B�"D����F*�5�f��;x� ��N<����d�&4�������M7��J3y���w�����o���{�g�."����J�܉����Q�)q�xa��>؄�.��R7C�+���*�nٕ5͖j�[;��-�x���ɳ�2ɷn'�����n�6��+�6_�l|iM�p�M��˾�|����e�[:������ �.���J��'N`5A��f-�T*X-�5݄f��൩@�A�t7
*o��Z�EG��Ne������(N�:�� ��[��[x�{��p\�ϟǟ���?�!"DX.�}=s��~�i��P(��ѣʰ��ַ�;�ۋ_��_d�P333��׿Ύy}���q������죏>��Z:�����,��~��y|���K/��ޝ;�����������_�y쨅��N'c8�����pxO�A6M-�H"uQ�L�ǒH��A���ж�Hv��(�]�!s�I��㺊d]����WӪ&N��̌�j�E�U߅/6�ո�ڹ�x?-�B�o:���H��H��C/呟9o��9̟{����f�6���u��~p/n;؋?��Y�q6�|qu�D���w���k��\눨5z��ScB/�����b��u�V<��Cضm[�q�<y�M��;V����Cwww�q;v�Y,fgg�H&����?��۷7%�����;�0V---���{��,@���7X��n��V��R'*��5M>O�L����<VDBD��4s�h� (��������_������O����3����C -ګ'�����>S?+h���m����~��Ur�M���W���ꅼ`���nO��;��W?��Y�t��A?4����Pc�.�\�A��$���0V#��ҍ���}�0�����+o��(,.t,̦=Z�'[�cqBY����vx�x������w���}�Ku8�FS�,m[����1�/ ;v���T�r1�������7�O��������#s�� OS��2t%X�rD���b*�;]G�}�Y���+�B�{zz�S?�S̲(��Po��lLk+�b�����ʜV��t��>�����h"��[�/�i$�d�y��WW�@{�V����ʨ��Z�!��D������ۿ�#G����n�L↱@�Og�1�WًڝoǛ��-�1����F��^�0�igw�1�k�]�0�����s����x�\j��B`Ƕ��_#�iMf�ҧ�VŊ���[>��}"�r��tY6cq�7]��;?�S,]~��8q�4����4���;�kwt���".�-���F=Z�0unW�e�Zc�+�ײsP��2o�+�f@EԂ��� �i�C\�fj����mܻw/���/29IJĭ�k���dD��LU��,�@�d��]����ge��M�-"jj b��u:��k��Ϊ}�g������D��0f�3!v=XA[�U�s���������7������=���w��YL���LĿ��P����I��0i����0���{�a�`��gp�|�RpF�aB-t���3���Wݻ��Z=��s�>a�M�{��7s�|D���:O3z�Ɵ�����8��ONN�irWG�yϞ=�ԧ>��~�ͲVb�8���5��m¯}tv��VYE��X�y��[{Ѷ�$;�i`�0����d���?��׿�H,8!6U-͂��}T�耋Ⱥ|E�Q��wގx[�+�bZŴ�%:ճ�������]���fJP4KB�&M���������3G��+D��F��bi�LD;k-dd�э	�aLsXA���X(J������j�A�E�T���ږ]+�_�7;!M��?��?b�Yh�����	I�Fu��I�V��ߏx�������6�$нI<|� ~�gvc�;�mh��8VV�'�?ݻ����LB�%�%Z�6t��?�E��;9M`Țਙ�YtX]��	��@2�ϵl>�D��q�Y��9G�C�����B�#,�B��?O����v���|�:�_�xO�6��� ����m�ţNra!8;E�-xT���ح�Ƃ����QZ�������"V�^Z�KS̍. �|�2���!B��uj�ȣ����U23Y}i?�Ҳ1���9
���żu|�`�r�k�yz�I/M�I>hѼ�k�J�Ł#�=)�X�܁M])����6O�evm ���ȥ��,�ܢKR�xK��ǂk��E<�{��Ͷ�Õp!>Aّ4�s,զ��x�h��Pz�n��&e��+����6������$�ď�`z��n\�x���wٔP#�Ι�R�&hA���0[H�H�AumdddY��F��fq��9Ffm�(��b�@֐.0KL��t��;�����-ozv��`���ʷ��m��6���j���"�|�4/�I��BϏ�z����23!�Z �E��5~i K�;��r��n/�@o�K���نǌ��N����MaI�������H�q�3G/�s떂�f�;�g�8�}_�^��
�|�X8���]�g1r>\�_3��'�4k��.������iF�H&�|`Ӛ�#���mJ�17m���oDMǨ���V4J'b��k�5L��\���c5@�&G�:��Ǝ�~����j���O<�DSK�S�^+��VJ;wG�H\4����A"M�6:�%�Oq�%ѡG��L��T�H�g��.��L=���\�M���m�G���,�.�k/�
��턝�,�����%�zh�Y)�P)̛a���M5��̿��g��Y�{cH߅k��y��y$d+��n�L��J)k\���� ��a��7�B.?�S;��i�{kӕ��	�߈z�:@"D��Ӌ�Ӱ�U�|n��;5"a�����_#�����r�AB9��(�|c�F�=XVc�-̡mr�b�z!wf��Vs���Nz�,Q�b�u<B���Q���d#azz�lA �`o�g>|�l�r�WlJ*7*��6�-�㤐P�����ҽ����jX��f.0�m�oWj��pw���BL��Q��)���g�[�j� u�<3#�_Ҥ��eɷ�X�q:�Ֆ�'������~p)�sԉ�vv�!�A����L,�n��գ���<��AM���Y�#2�y���g�y��7:ȸB��F����3�G��G�ڂ��tu ��	�Tz`��)�]Fn�Z6_�x�ٌĉ�ZQ�e�p��B�q�C7y��ή���.���_a�"Ks�g'bI���K�R\����G�G�M�ﰬ���3�p��3�R_}�r�����.,d��=����h�����kZ���j�4(M��r��l�u��&֔@w����[�lc�7�Z}���/�S�U�5,\x-��A�֛��
_�J9o��g���}#�J� �_\�g�t�W�f�9n����Q�2g�B�o/Z���t��(m�My̍3�mI	x: �I'�E�vZe�ߓ��ݻ�|_n$rq�L��r����]-?լ�Z���k*#D����fS[��j�aǚ�T2�{o܌��o;vln�ϲ$��� ��O��̱'�x� �7 �H)Òt#s��0����%��ÜeZ�.�p��[�,:z�Y��I��M��̑�v�Ǚ[;N�e�6�����܉�RXr���a�3\��ϑr�DŌ����=�X�w^G�u�W� [��=�aLw�2_�B��@��M��O�P�Չ!B�&:f������߿����7�����oc��Q���}� ���}7ڷ߆T�v�g2L✛<���?����l7��E�֍��SҪ�M� �ūݙ��i^���Bw쾇�9ٽ;�R�";v��h�{��qw\��f�$W�˲;W��<7Ξ�6|� �3�E<��4",a� y�O 1�Za��^�*󵀮����)�yD�V�	��f[�q��NF�\�X������	���j���MG� �$wHt ��4�h��J�l+l�${�܋-�y1`م�uLVmT��sEc�4gǎ�����5�Ci�����L�\�1�,\����y�i��|\�ҘL�[�잭��������` ȸ��<�2�4���{P-����]�t/G�����E�� VA��!B��Xu=Г��=���!��W�QW{ak)�4�[��hc�%D<�'L��D*Bj�a_8cvV�)��p:h�2�@�u�_g�����M�+���Nii
��)��?4Y����fa"�?ߦ�6������]�V��$_�+N��Tw]߇����0y�X�[�5����-��� �E��ُ(����N�X� +h�BT�"D0���%��)��Cho�n-�U��b��kǩl��2���M77�Zĸ*A�"Cu,uB�X���jlp�P��
�XA�|
��Ӭ4���l^n�Q�yÊCw鲝2���v�:�����F+	�̭��0��?=7�b9�Ե���c�5��f/,��,w�By��xP��r�6V�@Sphg'>���w�|�n��p��-A����&W9�*�Z��MHu�B�w'�][�h�e��x���� ˥\9����$�'Q�\F~���LB�D,��uC)Q*����I�f/�a͑�X~�'��>�s���ɉ�ݦ7��5�t_��p���zҡڭs-��Z@���$��Z�(�"DhV�@���;���6��Y��Q7�w�S�s���H[�7nI�e��6�X�-�עm�;�:x����)&!7s����mx̝N�9龲���#�\)1u9;üm,�����[S1c)���sT�:\�KV�HEtរ䮏�i�iO�m�&s��a��V�$"w5��A ���a��|�r���y�e!B��B���n;؋��=�D\�W��,;�]�pͮ :v��6b{6�a�}!��$Zz������|+�=?N��ihU��kђF�:3�p�Ǎ��w�����rcG1�i,�e;
����kM�f_#�4�|k��p��-*|�]x��<~��ړ�Մjёj�� �(����Z�%�mQX�2��^�A�_y��9���Ã*����1�x�V�B�w���߅�T�< X?��'�|s��[Vg�Y�&z���{ _��l�m[\]��-h"������u�zs�A�eb�7=/����2b�X��d+�ѹ�^�N3���-���N���/ϣ}+�U�"�bt���I]��1�b�$m���w���y�q6����.[jU�4h��B/�$ԓ栐"�4/G.����A�&�6��A�/^uC<��;B�k�'�=�	�U�5[�m3�h�ux��R��k8�نM��ε���HvBh<>��Y-т�-����O� E���ߵȳ�]>VE����=f���+���|�E��`�ߊ3�=y�2�~ٱDC�����X��Ű917���H��w]Ӎo���D��+�Lp�������Sϒh5ϯ%Q��4�5I�0BW���Y&�A�*=~�:h�a#aE	t<�ށ�޳��5�%�09'�n���68$O��Ǫ�q� �5��%�L��م����h��.v�oZ^�Tc˵BR8Z�8x��е�AL��wȎ��J��a��'���`�Vv�"�����t�B�T�Gn�+����#��H��ʴ�)����l?Gb>��_+�kMB��E�4����+]�9�[�4���-��&�[+���E&!�F�ގ��v��-)X?Mk���ZVQ�����粤
rH��������Z�nFP��OwX��w�G�ku��rW�,�݈���'f�3G��<yh(q��9[���	m��e!N�����b����P�V������8uy�7ЂB/�P-ks��_���4��u��E�e�%q��?�X�^��5����ea�����O�"Dpc�4�0xxO�i�d�t���o�ʰj�8�*�e�(sk� �p�9��H�t��=���_@��[.wn%5X^�׫�����T�����=�e@&�d'�C/.	Vb^<X�T�S�|%k�&\k���i���A�@?sd
�������ٯ%�:^/IR����zdTb��V�4�AN�_y*iG=�/k?+�<{���6:V�@w�'��w�^7 Z��2k8!�������!K�ݔ44�t�A��i��� ճ����QR�$?]��yW�jo/�Hz�~ly��`��/a��3(��H-k�.�TȦ�ّϸH6/oM���}�v�&�W�c2̵�FB=�� i�P�Tu,(��ǂ4B��4!�^��Gk]O�f&Dx�i� /+��'��D����":f�׷������ߚh��p��`�ZNh���ކ ��ܖ�xk/:�އ�>�|9�0�;�eXc�<V[�T�X�E�dKw���_2ҿsǿ�6dq$�'.�֮��#������̬Y�[��Y����6�[?���ƳB��qyu�AB-�IP�"AA$@"��m���1�D?B�&V�@��������&6,�l�1����.a.��hY��
��	j[^Er�O����s��m��[z|-B~ӕ~S��~�aU������H����G���o~Źa~�ɷ3���N\
�V��tFs~�6��6�#�35H�z��To��4Ԫ���t�^��zg���~3�sA+~i"��]+���:!B+B�i���
��uB4u�������M�]~�D�����	�6w_�0��#�"j����dË�֒��q��Ʒ1M�ѹ�>�.�So�
�� q�%N�хM���
� Z�]ؙm�/�K�!�k��w]�	���`b���:v�QK��w<h�O��N���UƱ�z���e�2>���5�0!B7�N�����}ۑHh�D��e����HwmE�s�T��RX@qa��K�K9;.]�[>g�g�&�l���C�/���J��U���-~֫���ֲZb�V�ﺋm>s�Q�\���m��V~�}p�f�W�{'�)�[��xn�=� bܬJ��ٖ�7����K�\�E�!�J#��?��>B��h:��9Њ;��e�2U�Z[-�d��wށ�-7#ݻ���#&W�Ρ0{KW^g���G�+*v����M�u�m�� �RN��k�����W&���^��BA�E��X��V��vt�~l��:JK�.K�y3�kM�˾��0��M�3�-����b�6T�xK��M������4�&*�y'j��7��\Ffi��5B3Ԫ��A�U�SU�Š� j�S��R�3r����j���i�5��y
Tm��9]_�n�F�	4m�L�Xq1���AC�g'z��:v݅�A���7��b��A���z�ͯ2�'t�},j3��薶@Ӝ�pL�O�}�m�l�c�N���X"�^R
/�G��
jN��E�����C��v�� �S�;�-��KL��5.��(��s��F�EK�A6����AH��zv�E���b���@�Y�l�k�������%�΀g=�VGT-�����A/W�R��:��{���|N`��� �jڗ��%B�����t?}ˀ����Y�i!_������raZ���R����dNd�x���>�0#��Ȫ�l�_���l���.5!W�A��IQ�����8����G�v�h�����j�͟b3���4���wv�G��f��sƘƽh����?[���bA�����B�wNyV�o~�YkԻx����j����2@�5���A�'^�@���a"D���h*�~Ǿn��oe�uK�L$.�H�e�zs�[��u�J�œ,���W���v�����L��5յ]�0���&)<^�}U1��\M���Y��������c�k�M$z~�ɓ�����3��:����w�c.��G���ۍ����ϜCa��ug�F�vvb��v�|zv��8�:ݰX���� r-;h?�P�{�V��v���[m� 5-xu[D�2J�)---���u�-^��t:��J�hJ�������2�T��)\V�X��[oA���f���ߥ˯�\X��%�A���Rmh��n����tQ�҆�O��XE�e�=�ر֫)������� �1���1{�͒qp������Bܶ�ϴ�,�� (ݷ������-���Mx�����à����k�.�R�����ynnAD�r"��ԴkZ���
A�5��M$��*�
�Ko��6VԦ��O�4n�����7����曈!��i��-�[��-�����p���'���'a#k�iA����Z:׺i:����>W�����X*k����d\�l���:��UY���%Ē���u'�S�1�#p�,3[��.��fTi��t�]��`��ϸ0�ތ���y�@��^�o�>|��@{{{C�PY���8v�V�����e˖���̙3x���199����� |�Atww7����}�Yd2���=��Cغuk�qQ����1
�Vd�$w��7L�)��r'N��j�����'?���(�T�W�@S]��S�{�o�S<v��y<��s�!��i�|?o�"K��y6��E�bI$�z���oz�\�iq�a�fM�mB�Y�ڷ����V\9~� �H�L"�UDX&���{i�e����^<��܂�]w0]�MVta�ai�gRX`�*_�x_63���,��ܼ�]�yn�`�om�gW���:::�w�^f��C-+(M��;w�	J3h����G��
�����<�͛77|^}��U#�4߬2����/�b�	t2�ĵ�^ˈ����x뭷V�@wvv��.}6J�ɓ'��k;T�c%)"lD4�@�q]�ɘ`(	���ס��"#�T�$�\� lA��⼏y� k�����w�؏�������U��\$�{��7P���K.k��r_)V��O��ܫ.t�cB*�����M�@�G}�Uw��X�H"������ŷ��jF�[[[W�`н��Ti���j��kh�ʻ޴/--5,�h~�i�4F�A���v�c����a$������6� �6ǪTa�Eqz��*u����̯4Y_��G�kY��d���Ӣ�f�«�W�!��n�v+�co�0s�"�B�Y�8����(^į�8�Jq	�f,�;��߹��Ơ�ʽ�>��<�����Y��U�r8��.�zPk*(y�p1�"��\ϻ���+W/C�|,B����h����I	�gK�a,ڀ#;z����>��x|��klG<��弜�la+:v��,��N����F�K��%��#�~$��ƻV��P�w����(�^d|�y�K.Xٖ�%�u�*K4}/g�Q��h�y�v����t��%�����A��L�yFke��P�1�sk�~/I�*���"������ ��@����/7�Z��=B�����vw�5���6�Q�e�8�"�0����Ւ0�ҝ9�UYQ���tڶfqz�U�ڦ�)�"���xN�^u�|M����|-�K��m�Fd���"I9\O����N�+zo�٪rQuB��K/!7u|
�AZS1V^x{�^��V]JG�e���}J��wC�����~���_����̛����@KNC=���Tm�@�iqn3ˎ��bff���"M!����D�A�%�%ZG~�f��#6��Y����EL�
�^�2�3�a�5!bn�NĹc�]����=�t`��Y'�)�W$~dX��5m�
+��+��|��a$��q�.<�L���h���}�A�r�'�9�s����.O����@?~_�����F@.�h��Zb93A!���9(���_�j_V�օ ��l�g�g��$B{��Y�r����/��_�r�qQ*��!��)���I��8�9�o��aJ4�A��E�HV��O0뱎������"#ϙ�߃^�����m;���$R�����c���8�Y�o�Aa�:V��r*��/����1o������q+t^��/z���wm[of2�*��^���ۘz�o���u�?�ˇ��{��^@����AV�BG~���abA�f����������g?˼P4
ZԶZ�&�'*�F]�q,..b������|�+̏p��:�ږP"���p���(�ވ�F�^4L�{;��ܝ2:<��r��P^�T9��ٷ����vۭ[D�t?T),bi�v>?}��me3��9K'�8�#����Su~��z���$C�����Za��L���-��8�,
�y�����5��q�D�t�y���isgBF�+(Ώ"s�i,�}�m�%=��H9���e�:���nӠ�03�1OLL l�tӔtA�d5\�5�fd��@����Sc!B�Рa�g�͒o8>��3�͏�ҋ2rǑ�-`#�Ķ�Z)l�m�4�3��hV ��u覺��,
�E��ɤ�Os�7�\˺�g��;&�w�e�~$�6�[o���n�i�ɔr�;�oȜ�w�YJ<�n<�<{&�~ж���ϟ�;=��	���ٕ�_!B�"D��Vh�@���j�6Pᰤʎn�$y�(͏CH�}�
����HumE�k�u����Ud�ւ>~�E6^2�4�aU�m1�W�Tr�4�H��Bv�(ʅE��Wf�8��La�yMq�R��#U��4�j�t�"D�aݢa����������&��!���SX�&2o�:~N ?G�ӛ�QJ)T�f9�J��5{cY�,�A/��u��bDU��o*'қ3���y82fWY�����<��L씹8:{�{������c!a�"D�!���	�P_�m�bQ9�r��ڑu�WVKlR)HB���G� �}{����:�11n/��Vv92�1�ŅrzŴ�Y��4{�~���1�vU�f!;��>�ț��(���߶�1�"D�!B�AF���;�d�ZD�����W�M�e�w8���e��,Щ�=���Z�d��x�ˮ��O��h��"^����'�Kv�Zο���7�?��Ɯ.P���`�'"�"D�!B����t,t�%��in�	�:'ـ�XP�5Ӛ�c$�a�c��A>eY����,�~8��E{���:/Y�� @eqW��K�x[Ӎ�Rr���������YqXR�aЬ�6��4ǍW�"D�!B��noI�E����դ�w�������X��>�3a��/��-T�����+����u*"/^�e�^��*�d� b�*���m�vd�j�@ �<-�eU�a0DA7w5�{8B�"D�!�h�@w�&�����z���g\��k���<W��KA�@'�7U�G��x����%�u�9�Y���3��W>丽d&�|����t��g ���p��u��XZ�F����m��!B�"DXoh�@�������!�����<g]�9$Y�N��o-�Dk�pNS~��U��T��1���g��%��n{šZ�X+�x�Ôp��sr�v!��^*v����7�|����*�!B�"DXoh�@���XL%X��$��9_�3t,ٮ$���W�Qk�_-�1?�]�gq�W:������c�N[�����=����ɲ��v>5�����!B�"�K4D��	���_{5��ۥ���P�WS�sY�cq�1��r�s�"�^q�Y�� �yRy���-~TI:�D���A��->/N�e�^c�Ӵ�m�#׆"D�!B��z�\�	�e���.M4��	�y�`��G���Hq��{,���
,��+��VZ����˫ul1�%�!����5�IV����]5� ���[�G�!B�"�G4D�+�jj��2$[�[΂�zL��̚� ��a�=񜟷U^�l!��p{�_���I����]"�v\�9�S�|3�~:1�"D�!�:ECZ$��"2pi��g�K�,�f<��J)_����D����#?�rbܲ���u������!��<P����t3^M�.j���\ �r%r�!B�"DX�h�@�*!TM���6���R���B6Ƕ㩠R��%�^�c9��Z�?�g=�Բ
�ZH���V�t،|�r��NU�ŋU�۪�����w��:��4��ގ� ��axx�ry��H$��ֆd2� �����
��+�����=�z�`+z�/_���̊߫���6mb�A =���yLLL��=c�`���T���"l4D����ci��Μ(;���󐉖�y�VP��� ����sL�C�E��,�2j-���ak�2�	���wLu��rnz��y��[yZ�/�3�����J��u�Vlٲ�ɠ�T*���;wnEI4�桡!���	N�O�>�|>�b�!�L�y�Ν�@�@S�iPw����ή�}(�;v�`�X�H$=sJ���؊އ?��A�?<�� �����>� >xY�{ѻ�����O��ʕ+��[iP��y�ftvv"�gOF��/ֵ�l=�1]��<��L��m�����VP�@�s�9y]΂B?�s-7r���,Ӫk崋�S-��y�ש�Q����K9����������*��8k`DBu"_\Y�+��m۶�� �g�mpp�}_)My&�@$��$I�k���N�Z�-ϻv�b�IP�N��ttt`�޽8{�슐h�3=w�cA���l�V�D�=(�t�kZ��>a%I4<i����˞;�(�t�={���� ��{j�V�D�F#*렀�8j����H$���w)��@���l�J�v��+e���7	��u[-xy���6{��֕a��k=��������^1	�,�����/{�uL�ú}f����@aܾ}{ �3��	�k�H4'd}��h#�d�Nn���M�DS�d}�4H�I���C+A�)�D�h�����NVQ"������75~ny޽{w���w������ɦ߃O������O�&�˄� ���L�I�����y�;O���'Obqq�����N��=z�A�?={j��D7�>r%���I2�jj��ԶJ�Y먎ra��	$��]�q�zk�����i-mr-�s�[&�����5p�ߴಔ��^�֤jvx��34{h��������_�0R#M� �D��!�}$'��I���$�����$��g�3h�D�s"9G&�A����u��X���"8�$�Kh��<����>�D�I�i�D� �VDP�)�+A�)���n���9hϞ���h�D7�DS}'�L�gz�A�?����F �����(�u$�	�ʪ��M�LkྈuA�!�v�V��l� ���a$;<�Z����V�O�[V�o��ZǼ��
����/fFl͸-��>���oq|#�5��:.*�ɹ�!�D�!�D�Q9�|C$�N���۷/����DSz�D6B�)>Z0G�S"��YDWW���FH4��=�-$u��h���Jx�'ԁ#��H^3I4S��ڒ�睓hj�Hތ8�=:p� �SA�?O���A��ݧA3����J+�K��wa@���D���N&�<	d��ܥ��d�K4�S�o߸Іc��P)P����m�8��\�[����˺[�4�+��%���^��4�.��_��h�\]sې�(�p��Ӆ��퀮xFgrh6�ӤF�wJa�Yy�r���s�)2j�c�p��Hy��FVc�ՒhN�<HɎ��H4Mm���-;�3Y��&p"�-�D$��*��3��<�$��N2������;��gކ�_.5!��«�;'��^{m`L��\��P[Mm^#�hny�w(��YD�������hb.�b�=�̙�O:n=�+@,�x��tm�X�����*�%�R�x�@� ;~��En�8[P(38�"]�'/r�"��q��,Ūkk�CNC-B/���@/����%��_⭽��s(g�Q1�%y?�-�|���2���Y4a%�"x�BeES�䩣^��<���>�G+��'�ԁ��<��$��/�,�����gD$�����0�g4��z𩩩eIj7�D�E�Ů�����e[#�F�Ep��A\��簐g�C=��r�h�G�4�3}�j)��΢X�u3�ҍ�m�Dׁ����:���/F��c�x��w�4�A�f�m^k+B*E�g��{��;�_�4�O�!�����Ma�ȯ߂B�E�}TǼ,��Y1��s����E��8�][ѵ��й�^���Y��Q6�w�⏐9��ӧ�t�Q��,�ැ%�|�ǛG��l�[���D��f�X�yM��3'�Ԡ�U���3�4�T�ij���3y( �$�yzz�.2�5�\�VP�9	"]/�����#y��C�%Ѥ'#y���=��;O$z9g"�tm��3������&�,#вE��o3g�41$;��s���>�3q6���d1�F��a����oa��?�8?j�o�(�����[H�Ǿ��g��V��N����+<�F���Q�W��f[N�W���@n�U�A���[vC��u�z�������+�CC���\�Z��̛_���g�'�U�8*�D��<��ب�Ԧ���N�9x~�>���'ܓG�d~�V)"�4��#�D��x���A��[�k�hN���=�X� ��?��"���k�z��dy���BK�9蝧u ��靯�DS;v��!�w�'��Q��4���+�����},��c�����ܷu��x��!fe�~�P�[o4ǒM�#;z��2�+��2��禍{����Z�?	��Zr�4���J+�,���Ik�[φO�H����]�C�{�����مޛ>�f	/�aSY^3�X��T���g�D�uB�9�Q�#5*�]����`p����E�����B�Dp��[��Ds�̽�'���X/"�g+���sI�T�E�����@�9���\�D�U��N�����D�Ex�<s��G����n���j7>N�M��-�an�� ���I�������X�������#��mF�����,��uO�~^R	�*K��J���>^zhx�'O�]m)�+�8���A��-\*K|� ۝{�Ga�<
�L�����q|x�a���eP]�4�Ds}�H�EWu�<s���K�.�H4�d4p���F!Z��CI4����=����gz�a�mx�d<<�*Md���_ou����7����PE�����B�9����E��ď�Ҭ'�W�0��:p��ޱ�mi��Ӝ�}Z�־�VČOٺiu�@��jC׾�"7~���Ә8�h�<�cq�'Hz����Q�j2��é��
_K*�W�ŁbZ��%dǎ"?sz�l�n��b�{�~^���6t6�c.����k�]p�Y��F��y��!��-�Ԩ��o&wm˅�#��qD��MR���`����N�y}���z$�"�D�i}N���z�A�$���"�|���u�$�hZP�u�|� �H������Ջ�j4I�l4
+�2?����u3h���%�T;Z��c�,��V�����U�4N�4f]]��:��ޏxk���zYh���-��^�ߵd*��'��mxi�i��ҕ7���x�+9ٱ��Y٪�ᕆX�ɮ��[����4�r��w]��z&�"x�B�(u(d��Ft=�#�@zp����G�x�"����>��b��V�@��@� �,��=�J@&�\��&�	���O���>��4pZ��C�HD�oD��l��d��x�g^�n�nJK}�|ټ��;n�4>��k�����u�~�D[�X�����S�K����ȫ�D�q�$���O��E���/����w�%�	G~��毘e��[�q6�0	[�YU�5,�왴t#�ha���{���\	o5`�&E�F �"�Q!�#}R�'�ԉ�68�%�8��������"����ݧ��2x"P�9i"�<��F<qM�
I9��z'�\�D��G�D*7�ш��0{�h��zal�m�1؛F�"k�uӏ����O=Ĵ�.,��I[z/^|���k�*NY��eiV�J�0�W/���^~�x?K��5�'�$��_f��g�����镲2U��2�\q��'./bv��G�D���U-PމH�Wݯ�� ��"(�D׻��4h���>����(䙃��&$�X��DMu`����#����lCͬ5���J:�<��������0y����HD7��_E<U����0�\�����,�"��i��}�9�%��:��_���#9�yI"�,�*}8�KN��j���K�^6������������#s��^r^UeBސDDP���?wl�s��64m���}����F�DР�N�<sP���y#>z�a74m����3��][В��`�5�L�Vҹ���:p���WN�y�E�e�ȏ�r�p���_�t�._����D>V+m2���eM��P�׊a���R~�l��������ĥO��-;v� �%�}�'���b+�%ȧ+�5����s�"D�aݣi��3���/����4���$�|6/�����w!�i�T�
\�� s�sip����ҡJ� �G�p�$�?�x����.YL���J�!�O���Hh=���I~U:�2�2&�$4��,��v<���N��8��3O��RTi�~&:��M~�����ܔŔӐ����"D�!B��;�F�gJx��,vlnA".I&*e�&N`�ķ�{�c��;]��$T/�0��7�c��� J�T�G����!ݷ�;���Z�� ��d��M�ȵ*�_|*9���G~�42��4w�����<3��	��]�ۉ�~�|`�o������L��x��?sd
�����>B�"D�ADSW-��kx��A�@W��J~�<�>���N�(� ���E��wQ)XM]p�l1C���,���av�d� R���^����^2	^$YEv��xi���JIX����mmn2[k�!�����8w�/��nz�;�`;:V�Y����c�}�	��������T���'��H�!B�"DX�h*�~��F�r�3����r�WZ�ĜA��Sg��*-�׳�������ǰx�EF˹y���&��*fܚC�`��.�¼q���QF��pj)�TY��%�*�5[)�I���u/�df��s��>��h���˪.�񙻻ɗ��(��};ҽ�K��m�i@�4�Q���0w���y��x{x��7*�ϩT[��Вn�{����'P,U!�ؾ���;�7g�R._���XX
�& -�z{Z��7o���B�R��"D��h*�^ȕ��k���vY���8'�Rn�y��M�dR-�6ϔ�4��s0�;����p8>>t�>LGia��٧y�:�~���
*i�9����Tq�hբI���u~2*30��g��e.b���/VH������6IA,��3�m��1�G�C3��2��l0}9��$�u����5���r01��3g�13�
�}K'n�~�A��k�B�LG���H��<[;�c[�^��pax�G��1�� ���݌=�6!�j|����<����%�
! �;��mK7��<�l���g&���#�hmI``3�o^?�Y����'�`����]]��)N��G�2F����d�h�:�N%�7�Q-.�19���h�F�O������	zoM踝#��\.�o���ɟ|½m�#�/���	d9;�ٷ���׹�=��&I�r����Be����xY|e��9V-LT�n��&����������gF�>����e.�P�\�/�Ԫ����#S���b���ّ2:�%twobV9G�c~Ve�4>'��0O��
Мvy��֖D\���+���Vl��û��BYh���|33#ZH�2:����Ņ��%�l+�����=6��n|.�
F2�b�Д��j��cWG9#��zY�*�y�<���Ϟ>���P�g-?��(���m�oǶ����H��b.N�I��=yܹ��0"�(�����Q6x��O���C8h佯��j��r�ώavf�����֚���N\wp�)3��F�O�1�?������sc�x��ߴt���E~5%Y�朸��8h1��k_f� v�1��-C&�"����껗����"ȵ�"U��Z�9��/�0s�8�7�qt�/xA#.��i���� �w(+�P���<���f�nT�M%4\�8�ݻ���CCu���e���K��2���"(���wll�P�A���Jļ�V@Q&%�ՕL&���XXȆ+�Fک����Fd04�����wI�����D��<�Κ�ׇe�D�dn���Qw��c�&6���a� �Ԥ2����4
����i��h�0e��۷��-+�<@����������1�(�f�7��nc�43���;7�?�^G$|z�,y^XXb-fH��,�R����Nk���v?�N.�r��3����9�\�KP32�ݙQ�w�2�}*���s��p��B��6☛�78G)4�~5�t]1(��0�{��6�*����Q�o��E��0n�iFʵ�D��^�+��I�o��I�t�b���.d����CN��%\��*�&S�0���a���0wx���Ѹ�M�_S8���݌:�ϱ����ݗ�1��V�D$ҩk��d)�:e��OO1�<�l6��B��|���^�2mk:ڄ�4���y�����yF�'1�:���|WI��3� �uK�ݡT�(���l�h��I���[�p��I�5�N\�8�=�7��lJl7t�XhBG;1I�y��_�-���x���_����}�^�,,^/���l���_4	$��Ig/L`ߞ$�*%�)����>x
Qۧ�i��%���3C
��.,��x�b����'09����Ex@$�����g�w��>�m���9�����".�L�@�X��C_;3���3�aw�=�aЄ��y7I��EJ�0��eҪ3y�؏����%t���q��Z�E\UVh�����u��?iK�1������e�[�4׈Q�<��"Q �� �[��t�`���n����r��dm�F��5������`]S�4mEH.g6"a#PD�h��K���c�f����$���a}���p���E���Tw�;��x�b�ה�eLLdy���F����c!87e�����Q�6OL��s�Y^��p>z��t���4�ص�$R���Azʤy?o�h�Ϧ�D�Z"u���r��H��玎g5�b!|�'�#i�wz�$�}��.��m�ʂ�l���q�O̲AXX�}��ߝ:=�����O�w�Ga���]4�}�</F��+B��
�����_�����ږ�6Qs>��t�LP�ƭ��F���̭gܔ�����i�>�ش0�6���|��%�����{�2�d#�}Ÿȝm3���E}����JH�.M�(�d�*�&�Uw6[��H�//�b"���*��lO����L�P�@}-�a �m-	�>3�d��H����1B�����^�E�R��gs%�ٗ���Z��y�5�-��u]��T0�}� �1��у��F_CkNd�����e�@M�d���5	w��Hz{K�O^���Ԭ�T�'&��`�X4ͅ5���h�mj*��1"�6�'�0C�ѱ&���F����n�iIW� �cssK�4�ť\��&��!�d�|��4�8�����Y�e�?��"jE��N���4G�c	�=I�4��e&���1��ߠ���w|
��A�d\ia�#�~r/wtb����5�F�g�|�o|l�.���p�<�}�ꆓ��+���/[9d}>>�"��:��U���#��7"����Q�4m^Cjpc��)L���l�3xk�Z[n|�m�k�����8�̦ќ���\�=��'�����q��Ε�d"�����@pq������p9��mIǙ�����x�y9k�L�����"�#o_��@s�����|�B	锰�8�+B�	�B��E�y=�ɘ��[we"�v���*�z�)jx�hD�rs�(\8��ٶߛo��Ѷ���1�C"�*���"@/�׊�sx�I�F.?{�?�K,���74�_ny�HS��;Q<�3 ��	c�t"�8�]�7~<�љM����Կ�����U��?�X[4�{Ʊ
C�t�v6���f��GQEc�{.K���I�����nÕ}��o�L�3��I�K�0��Z+��
˲8�-���y�v=�g���DZC�[߉j0�V�6d����3x�-�ȱٶ���#�:�S�U�#�cU�wGE{a�Y�����W���>�D�f��X�S�r^��Ȑ��~~��w����a[g��G��5~�"����k�9XVC��p�r�g��J"oYi=������'p�B�rx^,���1G:\�fVe/�$B�C�Q�Vu���X8�_Ϫ�oUgR�ۍ0��8����Bs�ܻ����j?�'뤁��[��͡X .K��;9��᠓g�.z�oZh���fI4�y��w>��
`����&�j0�T��}�޹�=�I��K)}��>sC�-Y�����	.qǩ1I��ѯc���.�c��H��AK���˂\�`�d�a�����;����Bv�8�f�jǝ���!�$ڲ,a��D�r$�K���1:��w_Ǖ��o&��O�Rv�M��3��uE̓h�q=w=}��'M29rw���0��ݚ]q��N;�9U��?dK�cg���B_!�!b4a��H%@|��50�&ۺ�_(�
,;��f���� q�U:;���7�k�`GGǊD^��8z~���{�6�h��dY�l9��O��
?��HCh5�Ѫځ��b��0�ɗ�_@���:t��lr�$k�U��ji��kݤZg���$��|��SX}z)/��e?L(|*
������ݹ��8s9n�өj�f�-���c8r>
�"4n��{bF���[���g��<w���XID�י���9q�7��w�H��i�c��b�;O[�9����1�T��OM�9 ���^�8+�}�W�B�q���]㵪v-\��l�\J����I\����V�@f�x���rMn��
OVi��芕@a�6/r���IH�]W�e/#7v�mN��ى��w�u�z$"�h�c:i�w*���o��YG��e�oǍ����ᗘg�Нy�g���.=�%��u���(�u�<��/����'11�"lk����9!}��ȺV�$'�bGR��)��
b"�	�����5&Ty��F@"��*���<x
7C��w�S�?ģ&�M��*Cu`=<pf�g�j��������4���nK��#,�@��������]��~x�ۣ{�ٖ�*��'���QM����V �r����zq!��RB~���w���D��uH��bD���[�c2�jy���(:*�*�y�sfm.�#?y��u&+8�t�JXF$��pi���5���o�����i�u{`�:eJ[v������ZX�I��3�+���8��&�������:��k΋.�	�"Q믓qf�Πj�.Z/B���6�(꽧�I�6�Ｋ�s���B��Û��@݆��q�H몺�A��"A���
��]�v��M�k�3G&�}�x�]斘���0����t�1���}ܞ%��}/�cs�$\��Ho)7���c�ҋ������j�mC��L�mB,�a��m�b	 ��Z/3	-$�r���H3���f���S<'v��~��ba ���r%��A�7���Q�s	�2S�+؜���2�p��n<�)�n�x����X"���X�w&��A�G�u�0��Z�-@���E�܎Ytepo�]��0��B^j�Ja�l���N��}�;���6��X#\�'�HB
�/u[}�M2ן�ߴ<�j^���5�`�9E-	i��ZH��k��f�o42���ύ`�P�����v='�̙�[M��6 ���K�(��	�p[��rn� ԳȎ3��X
�t�NS+O��/��@[�V�KL�L��E�k��!$"k/��(�6�
�]�--�����P��}|�Ա_��"�'�݆X����O9�K!��J�8�c�'V%��a���xH��Q7�v��P�7�b{����X���Ǭ\Wc��f7��|G4����h�ę��u;�y�ʊ�7 A:oCl+C��Wɒ�5R����^[W-AS�N�M����Y�ZP���W0НFO�t�4@TN-k���Sv��e_e$���Ѷ�Dl�l«��=1X����\`�e�si \���Uc�ҹO�2��4'R�FR�!_�ݐ���g�"�Ӝ�mM6��>����6ڑ��n���a�?�#2�F$LN�ulR,V�JđbN��ېD���T��JE!-
#�i|j�����X�yI��#��ޚ2g��w.,���teL��'ê�u$1$�g�n�M��'XR���Z'�c���<��/ɖ*�'o�wQ}��ٳ΂��4V�D�߆����E~OvNV۷o7	����W�5�|���>�=�m���[і�W=�h	�5V��8���_�Il܌&�T�N�B�{�.F�˹9�g�bi�uT���pY��K�C��W��<����"���"�m�Ԑ�����$��:�.��<u�F0��v��J���؊W���iv�����k��S�M���&�+������J����l���4����%�D����
�E[�*���4��^x>Y���,ff猁Q}�9�L�^;:�ӌL���g������g3u��o�hoALk5�!�G�Iڞ{n~	s��}�T1�3�~�"��0��������늲��t*a<�$BO�t�0/f��,.�N�>��6��"#�y�k�X1��L]9!�Q�x�ө��B��8|���z``�Y��;��7�2��?����Zp�M�Y��@i%�3����N�H��4�Ւ-��y:�܋t�A��tʦ��"
�Wж�2'���9�ӽ�z�.riGv��;�����*�I��&ZXz;v߃��� ��k�%�w1s����8u�%Cqvs��u>}��>h�'�u?99Þ�~=�l��%\����,hK��ub��\� @_O;Z�!%Ѥ�/�,�S�s��HD����L�Pbu��%Z#Y�G�f��i��Z{G�w�T*av~��QG�h��ڞxxd�3s��U��Y�c�E��:m�:P^��_�B��9�=�"�.�F~��V'�!����..pyt�<g�a�v��%��f�����tha���Hu?_�f���|�X2�@Eo3�y��8�����/Oar�x�+�w=��-i2Y��ڑ�⮻�2	4Y���U!��,N]^�W�����ޱ�ۥ_�s8�G�A��Y5lG`��%���{?z��0R=;ͅ~"�ߩ�HunA�c ����q���&Zp���6�d]��:�Vo��1�I����s�CH��bN��:�x
��=�\�}3�����v����@�:bM_�S��E_�j�xɎ_Z����N��Ԉp�l�xQ�o������y�D�E����aҜ�����,��^(05��M���6P}�26���i�����:R���`��i�"6���:Щ��9y-��*���+�K�@w��l��Ҡ�id���J�<iU�ۙ��xީ����'�=1�V����&13�q��ː�U�l���nC*Nm��\�2�ڱ�vNl��w�X*bfnў���p���m�Pf3��h�W����ο	��߅~�u@e{���^8R�c����*7/�t�tr��Ֆ��-��!�97�u�Dnm}o:��1t|8���i`ۖw��,ƞ�CT��V�r럹���_�$�獳���lM�&�߾�V�f��!��f!4gq�ѣ��Hq�/�[}����J��e���V��v�.Ld�/�g�ST(�yjfdy4��Ŗ��dvY:$:�$�����a[�\S��wH��M}+�3~%@�����{Q�>	����7�n��{�d�<mg�������Y�I7N�H���(�W�gy�gȠW�y7���Yy��/��]!@ds��ix�s��>�]�FN�h�X̚��t��p���D�x����yϢ�d�B�I�ef�4 ��p�L��ӳ�w_�}R/����ݦ�p����\�o�>�M:�[n��6m���Ԫ$`)_�SoL��+�O?�C�-�[:ᶐZ!�e�ց<c���}.+�����;�D��wa3t�D�����Y��!t�,'��K,`�&��B������n_,V��J�hA��h��.̟~�1�%�������l�Y��z}�B�VAi]�_�d�~�ԭ^�x\7�$YeJ����i}��/�B��1@I�\�WF����Z0��Xc�G��C/��ׯaՕ�m�L�ޟ,�K�,#��A]h�9�YD�� ��|��48��Y5�I_��Al�˕���,Z�p����R� ���T˳�.�e���R1\���y��O3	���z4c����Qoh͈��Zo�X"�l��~�ٝUe���Lc&�詹��V<� Z[[���lhh��?�����Z"�KLc���c�l�&�L�H6�����މt�^���F/��x��u��S�3Ӡ���[~��G�B���峄ܱ?��R�c�������D��m���|���l�­�U%f�Kl(yP��Y,����_�gB>��E�!!ˣ�浀�'F����Y�7� �zV� 4��2Nҋf���rH��NOg1;�۲��Q6ڎRh���˳VzKR��&�e,�捿J($��|�'�/�]�n&<F̞���a���@���Lr�|��Odtlb�8�M���=�Fˁ��@�lqe��G�H$L	����>��h�pGr��t��1������V��2ɶ��'i�i�@��kT��NV�D� �^3��
'�K��W�{�6�<�s�;R�!���j��y���D{?��.櫺�~b<��Y|��0��}j���<�ZVi�{�V��\U��W=��\�mTW��OyNLf�\d�hKV�syd2$[Л���rhO����Bob�˨��?cq��æѨyϾ��ɷV
�_=n��f��^@	� m�r�ԩUM��\_��y���"�m�h]��W�%�K�@K�k�Dˮ�=�D<��h�H���u]���A3~38�]�L��7���j���.W��,��H4]khY.�������T6_�7����:�����Gt��6��������O���<��Z�эF+�}�C���2U �$�d������~�E$�O�����w��u��~9=�����[����1ʪ��NdJ�s����)�:Lɉn��6�w��c;��qV���b�����^`-h�9���V(����#��>����cy�!B�"Dhzzz�?��L�L`,��3:��#���_�2���W=q��E���g����;��$ڶ�:��kC8~��8�rvz�V�yIG�޶���⸽A�ＷKӡ8���	\����RX ��]i��?m���8��ҌpOu:��4kL+��O㏿yn],�!B�"DX	|�d88�Jp"�I�={�������&	�dK�o_;�t�䝃�ܙ��9��H�{9E~�,�����C$�2yf���X��c��͵� ��7�����u�lC0��:�ȥ8�r��v��Hsii
K�o�/��=)�,ۀmY�����Y��v!4��"D�!B��Fww7>��O�O�*�D?[L����ܹs�{���u��wl�;c�6�pui�"@�FTJ"EI�BPB�TiՏ�ҪJ?��D-ME$HS	�&!��$� &`b��������׷�v���Μ9�k��]{fwi���zv���s~�缇�CC� 9YO�:��~*�J�����D$���%�/���%�d Y7b���[�X�Y��\~^��`��6���evV����S���āTv��Y=f,���^KކsF�bM>6
�����������}��\�G�--�ڊg��T�{��s�ʕ+�
}Ҿ}�D���2�h���EYUUU��~z�7hp0~/q���ϛ��n�f�rZT�'�����Đ� k�i����+���.���"-Gu��@W�_�3��&G�!��� �w�X(�htPj% �m<��|��b�XiP^�E�!��u^~O?f_h�d�p���Ab4����ޫ�onv�݄��|��Q(/R!�=&�������~���T�\.;�?�"�S�!��`-��;xJ;���t����S��\cϞ=b���Z<��^�m۶ѧ�~JgΜ��B~u����2���+h���� 74��k�aD��#�}��4g�.ʞUAZV�HW'`xd�F�D��7����&���K�?͒k� v�=�J[�ls�d������:@u^�'�=4{���#���)0�%�U����h���ø,����̯���������:jh�e*���.jjj��
�~:4�� ǆ�Е��TXXh�rS]<xhoo���^a!�;wnZ�$�#曠���ϧ��R�Z��}��G������g����s��#6-� ����)��4��1��=�����o��hc�E<( uT��4�V�XA�?�<���PKKM���t�OW�������h�lsmz-bF����c�߹B�S^�*�����P_�E�����2� &s�D�� l�K��Ʋ��~dG�5a'��~D��T�h#����2�犬"�:0�5}C��K�c�?�8V`GԹ�{�NV��_�ܦ�^{��kmm����=�������)��x�b��=�!������t��=Q���:Z�dI�C4ʎ;.0���`�Cy�͛���X&ZG�����✤C�!����<���SYYeggS:������Hb���]F�@4����&�EEE�`�J��Qcc����,j�q�!u$����~�V�֭[���ȑ#":4�������:�i졽�Z@K�� Y:�hŁ�^�i�}w�s�C��/*�"�Q밺T7�1�(r�ԥJ��+[N����~s��V��u?��u�P>fs��9:��(7~�c�4��5"߳����F�����{<���^+@���.@"���ݻ�r� �T�h�'D^�!�\{��T�H2<�����" 2S8�G� Q(;@J�fx��	��ǭ[�D���R������Cۇ6�Ν;�������A#�g�߳�V�\IA-H��&�@��MZC^hd���*'O�_��VA���mt]��=[��U�T67��23L�%/�E2�j��xJ��~!�!�e���z!["��{����Tr�
�Z����<��>���8f�5�D�������A��6S]����� ������R�
�3G^�F�!�#њ�z �� �� !K�h�s�t����������l�H%1<��3<�Px ���!��t�h��8��=��h���q����.?"ѩ�߱����&|a�ذa�h�Ux��D�����l�K/�$.puuuDg7������ooy����E�h���I��pD�{f�;�j���H��k�>˒�V���5&���I��8kD��w����CV��ٚ�q��( yѨ�����t�F��R��ɷ�RA� @� ��!D�����m�yV��XA�d*H��X�'�h��T@0<s�W�?C4�WQQ!���R2<��'H�h-� R�g���R��ug���;R��ر�b�P�l�$B?��{˖-t��!��]�r�#�?@�tH������+�_������+Z��hV�@�"�&��%k�̾��F���e��A?��mB�f|�u��	��o�0�l�
h>}�(质s4��-��9Y2<��8V#��s8]��3��r:D3<�>c+��jip:H2<��֭\v��8]2<�6x�y�E�pK�
bxF��ȳ*@�}��+U �m>�4xf1D��T����{�- 3R9c ������%����ܾ}��>|�jkkm�~���槣�oӅ�n�՚�Ŋ"Z|_�f�������:P�����#��c��B5�o�]�}h���<�Ȉv��B�l�#�����U���~�N5��404��D�#�N�hnD�g"��P��f�:�h��X��pD���đ=^xf1H��Ω ��<�]Yr������-�!}G��,�y��hB]�w�O�H4�3�<��䠑�!z���t����{�1z��WE:�Xl<�Z~?F쩧����o�- z�&,C}��n��쥯�wҦ�bZ�t��h���iz�<aϰ�&u&럚v��&M�S&#Z�R�)O�mm��5�[4�:$��7����:�J}��4��Byyb�!z��"6�7��ȫ 9E2<��8��4�V�y��Hp�0�r��A��2�>e�uw� B�g�a�����O��q��g���/<C(�j�p��~O�(nW!}죏>J���:�Y�F<kh�-C�X���{�nqA�z�-���N'��o����`���-�Ck�̡�if^��eCS(lT���[�pjP(l���/��3Ø ȓٞ�I��N>�d��(�E�����C��<bЀ�N�9�+4��P9;���F9�U�/<�8c	��|�N����3�ӝ1H:����8���rDs�ǵ<��V��?�D�fx�ǶM�Z� ʉ���֡���7]�,�yuD�]�)��>.��^{�z�!���rY�\HE�h�h�Ry�gD���7ߤK�.M�SL�<�a:�]']�A���j�L���i�����'��YM4G�C3"��DK��l��ߥ	��mC���Eه������m��.��hF���!i�%4��2r�$߷��l�iD�/�At���x�0��y�t�<LvEW�� 9�9�e�h,f�;�'j�Q+C��<���i2��8W4�$��uC��w�a"��FN��*ól�����O��/�L>��ѯDK��2,L�*D����{ �9v��%"�G��S�N��n7�ҀL�t�<w��(˧fҚųhU�,**7F@��Ca�<�/�ђmC2x�KZ-"���R�}��r�����A�ϵ���۽tY\k��;>j�����U�2����]!����F��'<���)lW��LĶKN�ht���g�$�
�܁&2]�� iw�V�|O���.�-}'@4��<ߓ���g Ѹ^ G�S�](���	-���9��m�	�s�^x�z��gE�T�n���Ȋ�ꛣ8.$Z���;��ҎҁY)�a��'%�TQ�K�*
u��I+u�.��ݰa\��|�2���D�4K0hZ7Ԥ���iTF4�	���40��f� �{~�u�UHhT��kv���I�� ��v�Ds��h"��͞ZȎ���Hxf���ގ ���[����\�2�B4�}\�hy�'*������C"�YާS m=�}"�����	-��ϰC�[�Nd��"
��e�͊Hc'�8�ӲЀa�o��ի��wߥӧO�:dZ��+6���9�T2;��+�@����*K���s)gF�	�����C�u�)��	����?�֮�o���� ����R�g@@s�ƚG�]�> �u�
��9��D�����o�hD9�eG�f�*�D�3ˮ �h2���9D��@'��ȖȎ-������<���n"��;;��Kf�(тs�瞣�{�
nŹ�������#K�h �>����'�|R�G>��#�����Lc����L��tЬ�b���4�8�*J�(�ų���0[=3��!�&��U`q���!���7�q��Un��.�P�8��`2�P�E�xō
F�Xz�.Bǉ(q2��0D��h�<�l3�'��d?�������y�煰���. � �z�̺/C42��i��k��ȳ*�B4��~.��,�]!����D�3��;����.�%Bh'y��]�v�����FK�˅aY�P}1Z�Y�GY���#���ƍ�ĉt��1��nw\;z��e����Τ���Ɩ��A3�B�r�D����t�́J([�O���m(0B���6���{����{���I	�
��.�h��l2�v �f�hөhD�Ӗ��M'��ܡ�E��SQ��c����O�&ɾu���Kf.;�)��'�h�Q����{<���E�[N��ϵQ�瞞��3���W^�͛7�I�����6��@��5�P�h:�يX�a����t�R������bsBDZ����cd�@ Z�Ԙ��e��<���)�]r�O�PGs�|�k�� �ɲ��](7燷���.�]�dEz'��*? �`�����$ܕݴi������SyyyԤ�\���ޓ�cY;b=V	>d	 H�߿�������ߧ�>�L� ������:#�+W�\���Z�R�<xL�k?�*++iǎb��˗�,�����9��h�#,*�f�%�p{��!l�s�N�>w��={�Ο?/f�����+W�\�r�����5IV�ZE[�lg��C��d<��ZPP��e�ɢ�tĒ|��o� �ׂ�^�}���6���͛7���<�QjL��1w��ʕ+W�\�r�^#����	��-[�Ll`ɪ�*e�e�B��fԐ+M]����0=��{��@    IEND�B`�PK
     �J�Z^R�#  �#  /   images/e96e51a4-2e0a-4cc5-ba63-cf190e1d4d54.png�PNG

   IHDR   d   S   i��A   	pHYs  �  ��+  #XIDATx��]	xT��~��If��$�d�7�b�\P\�֪�j���j�ť�Zk�n�Xp��� U�M@�@X$��}�5��L����Lv�_�繙ɝs��}�|�9�� ļy�b�
���B����hA�ňF�eV�6����U		�ԩS���g�}��g䟵k�b���())�y����5-	#�ci�!hj��>^��K���e�
"���ݎ5k�����/��;����|��g?�!Wē7e�s�"~��8��}4��'V�AhBl\.��Q\0s'�]��[|�sk�#t��0 �?�����������7���d#q�!����Bm�vB�nr��ap>\����
��{^��w�*�#tH�����0�Z��{3�lğ����p4�\��֊\8��#<u�Ih���^��c��\�p��a��;���g�!���m`�X����fq*?�9l6�)���͛a,//�޸�¾�ߌF�A�F���bU��r���y˹�U���/T�zO�0�.$E_��9��鎄���.�Bn�޽^D���EEE��h4"**Z|��Hݯ_�kc#�m�^�D�%�\�9s��؄�;wbٲe�y��>��HOO�
��7���I��l����=K0�����(#��`�'��GC�6D���~LPs�ߎ��4�yưD��ǯ���ǰ3�.`����ǘ1c�r��a�TTT$F᭷�BLL���*;vL"������<)k��'��w7c�䡸��W�����;���ݻ7�M�&K��?�=%22�����`��Ѓ�c���ض}�Ў�##c~��_�2�	�w�Fw�K���E��HD�~5�A!�WC�仡'������Mp;3�j�CM8w�gm$%%�{����<	����#<<ܫr)�8k:
��س�n�L@I����}+�~�J���֖�K�,����%A�nBB��M^,����*++�>��o�B��蠇5��И��(G�Qt���ƢL~���p6���v+�z
V=*�k�؏Q������ٳ����hqq��WSS�[n�E~>|�damԨQ��o~#	��SO���2`�M.'��r��=���|

�\Zhhh��l�!(���+�ȾTUUa�ر��͕��V���?=�ج�(�˔mZ�m�$)��Ê�C��r��0�C�D��5�&�K���eF�)6G���\ڔ$HPP��G�� ���/~!�G��-�P&�Nr7��hJz�[J��v�O$����7ɲ�bY���n��$�^��ֺ�b�s��X�,��d
��Eh�d��+�@��m��!c�B�ɀ��q�(�C�Ŵ�.2�o�\���NO?�t�x��;g��-[|d��I�U��S����>�*�T���l�@r�@ɲ̖q�{��� �U�B8�#i�ը9"���R����<C�4}.ly�P��>�� <W^y�do���?��,��>}����F*�C�9r_�u�cwYp��tI�FW���y{�k�m�ڣ��ʯ�7JV間*HN��N;M������;�q�ij�$�ɒS�9R�2��$�e�;�%��#�MF�Y�nٶ�#~�-���6+�ڿ\�ı�g�j��E��,Oyq��!�&�zKP����W�3�O����(�㙧�{���9G��,&N���lW�!\�?���%{�J�����>�>|w�yz
����@-��'棾� ���;��e������:{�r׊bF�7�a/ۏ�wW�� ����@�\s�5)��I,�&�2�
�6����[�n�������)�����Gq���]�P�5��F`%'͑�G����Y�r�������o�vo6��t'8#8��$"@\\&L��&q;
Ja��k~��gGqƈd�	���2%���?&�?�t���&�Fhl��S`�>�р��&,X���=_~�e����)�
~%������rZ��,��ʇ �v�}m^�o���6���z/J�e���u.Z�G"���(<��o�����{�7��C"sѢE��o$B���{�^��*#�ڢB�"�Mń,���u��N��s곕��:Z��_؉?�<S�w�>{�t���	J�6�YW�ڽ�Y�y�V�[r���Cj^�/�#�<"-��G�JWDD�:�,�8q�v풬���v̬Y���G`ҤI�ߐ�i�"--M����/e�C��_&;��/�ĬiŸj�v��pK��1��`�
�a��bk)��)�+�
Դhy�����/�S%��O��NK��"q>���s�9HJJ³�>+g�O~��"ڴin����
��I���ȗ]v�dCK���E��~�,�3���B~�G
�e8�����֡� ���3��ȦMEw����ɒ�1���oJ[���ߗ�3�[$5�w�yG�A^x!^|�E���ŵ��;]nd�ɫ��NsV�#��ղ�ǋ---��u`�)3��;v�{C��n�z�I$����?���$"�J��̙3q�gJ�w�ʕR��s,�x:	��������'i��߿_�"Ύ��{O:�(����=v�q�yz5�K|��ɲ���D�8�º

� }� ��c��FΑCr�|��dgg#''G��ʶh�q�N����^j-��I��lĈ>��ٚ�Nw?/~6l��8�믿A��_5�e�9�P�]~��r5�$@�Eb�����(5ПNN�38Db�b�w�y��g�ҥ�͢��[/Ù��a�Ɲx��%�l$aX��*��d��=���:�ޠ� �W}50����x��"#�u�N�&w��^ݞ8z8��Yp�b����^+;M�Hީ�ҫW/���"X�����D��fҪfV�8}_Zؽa!�O ;��J
H�sT�����/ȶH�� �j����a��w_$ң�
����e�(0��X�nK�D9Im�MY�\
��~��I�o��b�.m�ʿ���i���;����{����Bttf�5�HƉ�xD�[���!F�>ԃ+�c��O-��K�����-1\Y�o��7�}ݜ��w(��e�~���o�{W�j�aŪu����K��6�,fL?�gv	��bM=GjW\q��tg������O?-�r����Իo��V��w
Of��۷O����ӧ�O�ɵ6�L�<��CX��?�2@YF��5��+�Hb��u�qXV^��W��s/�oo���"���T�?+RF��/�#g#�X�
�&xM�nʔ)��㏥[���f��zh8X��&A�h-|��2:Q\\(�'��*��$|^��{��
1�ٖ �P��K��#�ZVL�i�Q~�\�����T�[�e��M�Fr����v�@=���~�oڴ�UY�F$>W��D|�[L�&�Ǎ�Z`�a�*+��n�����M<��XY1�X�z� ���Ѿ�=�6o<2��G��}��C���w-�����Bmh '� �)PZ��9��(0��w.��l�*���Juw:]�`l7!A��� �"��[����%HZ�t�{�.lY�k�<���FL�k����}����H�t�9�T�V�#1�hl�"<L��T$b�%�c�ܘyAo�m�^�E�1�m�GPp�%]__/�qv�=@mK�#��9g^g2H��rH��X'ggG�"��l��fd��=��%Eƀ�9�3M���¸�B/.ǥ��_�/ƺ�zX�B9	�F�ѻ L������M�I�"�'��м\-m�N2O�7B$s���̜*=A.��b����O��C㮻��_|!/�VFF�7߶-`{L�ӆ�+�˰�Oqdw��Vב��ؗ�X�rV����B�	}Pj�([����7�,��Ҡ���Y��)�)����}��&4�L�{b��o���?E��R����W]VxG��r��%x����1��m�.���t�y��Ȟ^�p5:NHO�Y+�D�9į��q���S)9����@��z��D���G��bG��1�|�-�l\�ՊeQeV��=�ba�V�Vnr�y �?M�C@aC@���A�+
Q^T(>[��/kğ�Ob�s��NQ����J63~�x#�"��mΖ\B0[,a����>��r��% ���KMMä�8vp�\�\�i��Ď]y�M�m������g����9Q��/�qm=��	r�D��a���=�����R�!-#N&�y�APcbx�.=�H���Lof��A�q�ݳ�n�j��N-hڥ��/�nE��N-�bڪ�!��n�q���Ͱ���sd��PC�����%HLL4���:|��'y�;�ԇ��#���C�À�ޓ���i=R�u�(�DE�g� 	RZV�vGAg��Te�z+��D��E׏vlj��0t��%筎�����"��S�
D�W�w-��bn-�}N�g?E��zk��B!��f���sʺ�.�H�jl�s��lv�K덩�=/�,S�w/A


��Gި@i@�������$joQ�i4���K�T�ŉꫤ;����k��T���qlfN0n��=s�a��O�ÿ���=�eYS.����Z�5k|��'�9���ʬ��l|��i�2N�믿�Sx������%��wl���>��-�l���Dl$�B=>.!�[ٴ�]5�3��,�Q�ׯ�j<���)�ײ^r�Fc��ab����B]�#*��$1�e@�Sg]2������D���:����+�>�����9�|t��[�[��*1�@�`�g��LUB�Y�L��'V�6ZSS+��`1���I ���H��>�Mض�/�	�ei�=
s�&��j;��P�>K���@^Z�����]_�+D�D`�P�,�o�ѳԨ3ڨײ<ĕ=DOB���YM����>60�ʎ����eU Я�1v�b��ڥD�*=�*;���	E�v��Ro�=C��M7�$�!��c��IvZ�;�@7YV��	�4�A��jY,u"Hmn��[�õ�s�N�d�NF�*�D����R��
A��!��.^�D���͌��ɨ]UL!�R�$��� ��eu�R����b�h�چe߾��+�y4�(�[���K��g����#�����O���g�׸=��<�Z����g����i�����l��9��	������X������\YD�rQ0��i8z�p�ق��4f�k5~gnnGd�2ִ�?} ��w��z@hq¢c��z�~��o=�-�=�W��,����[�,���͉�Q\N���dee����nj��YyT���e�2�'&h�D��i<T(���� ���Rc��N��(;f̘!��,�g�y�GYQħ��CjY��
�\�n?ܭ���@�׿�U�"�Lz��G����;P^V��/�Gv�=S����}��c��t� L�&��r�Y���-��ڠ!۳ګ��$l�Lz"�!�>c��X�J������֓�,�(�� �������|�,�Z�����*�	d&�>�K�%���Lv�P=MJ�PQ���u��APn�[����i�3�&:�"�'+��=���YN�A ��� �N��_=	�!��]w������L�>����<�3��� �:��o��� ���o����2�F[�[��'�j���J�ࣼ�o&A{BPG!$4�y�
���؍���<����\�#����e�0�-�qi��o���e�m�P���n�%�'H��gEG��H�?���TI��qE�=J�W˲��"g�N[�����o+���^�������&
Wjq*4�{��֙�i'x�M���@�2�(9�jW�j�&�̲TF�y��T
)Ə���L!G�<�� �w.�-))}�h�;�ڋ��/�Jh1�O$�'�ͭƧ
��̸��B��1�7II	2E�Ռ�℔+�Z���$^/�?"��� u��Ґ"����
�>���<����N��F��מ�9�;��;��0��\��R�>�|�X������A�]�2��[�I�RO����gi�J���r�촷���!��j�X��"]=-���b�����ib��w�Z��ʪp�sd@�Z�l4�hӧ[�n��Ȩ��'�%�;	@��'�Ӊ¢�n��� ���6l�7z��kq��7I�6N����8������_�~(��m��*��H��
�vyJ������+��
	Ow�Ί�w� }���oF�� �:)���WV��3�8C�1�����=�&�ic@	�͌�LH�UӒ0�,��C����m�c��J,�X��[��p���8ՠ��w$��$յ\*~�N�ւ_��	|]Ź3�B��W�x�"X�s�t��46!W^:�_��W-�o�y��?��6�}��'�2<�U�z<�����Un���Sv4<���?n
��楗^��q�h�R��.l�����񫯾��?�)n��V�l������ Ƅx��G��)�#�<HA+�K��'ʥ�#8a�|]�)g#��ʃ���*"�a�7C"mB����X�yyvn�j����g�>��NR�Q�����BrV��jd4NY�V��m�g�?����rP]և��vg�3�_�GW�)E�f0�ǶI�m۶�3Y�Q���C����x�p�&X䙋�}��P���|D��cx\�Z�*s����p���
F���b���6U�-��1�F����[�YFK�����Z`]�̒PZ�L
L"W#�H�ë�ND�힌�[�N^��{Y��F�AB_v6V��{��x�1i�rΆ
T�~��<L8H��N�O��+�㡷�.�6��ˏR'<�|�ٽ�4�@Ϩ��ym]�m�2���:�%HZb(f�7
�㯅;��h,Β�#'M�U����k�� $*%����W���xc�1d�?�^�%Q����@Hj/���}�O6��2��c���z������'�G#e�8D�N�`�<��٥�q�6m�-������0�F��LM��1rE@��Cˍ�0�-[
x� ��~�?��������s��v��kUD2I�LyA��bu<H�J�Xx��:�IE����z�"?����e�d]=%�;��U$���&4X�DC�V��`�k��wM�?�(f�L}���u�Y�� |���8�>��_��Gɽ��ZΘ�O<!�k7d��Ƀ(�D�P�5$	���
P�D��o��rGm��O�� �b�B`ף���$��h���� l�o١*\sh���$�X���z �eR5��j#
[�h����oR �iP$V�]ç|#�>��h�`l-����f�f-�#a��]�&Uh�ı�
���L4�nIc��TZ����}�
Q���f�7�8IԪ`_yԔ�Tj�N�_ڪ�v�mn��v��/Aʪub�\������*"�ϔ�֞�&ѯa_T��;�&�	[�*�gn��Wg���(Љy<����ԫ��|R�R����o+c�4��X� "S_��1G�9r�"�e����XF����11�e,Kן��.4�#p<���W5N�.A�����G��
y�;_C7�B�e*��ò��V���b�s�:���\�gL^�JsSs�28ؓh�YF�L��s�e�S�`�hN$���^���8Y�p�̐�
c��&�q$(c[Ww�7LͶ�H�0��h�w��IT0H�0���ғ��j������L,Õξz8��ny��l���Sp��m�VY�����*�j}Q�E(��
��|HNY��r�2��o+$�B��f��,����J�WB8&�K�	b{��pn�̠W���}S�1bhoI�̬����䲗��2�O�!��/��ƭGQYe�e8��ʘ86)�cPU݀M[���"��1
�L��Q���!sO�|��/M��`̈>bŘp���r��}zԘ���d���#�8^X-�ĉ�)�Fj�h�(��q�U4��I[��ղ:\Ԁ/6�bvp����F�\%Ά2$N��q�9�_��.��}�yߡ����X��{�y|Z-/i�i&�F�r2��֙��$BLT(�C$��!�>eTE1����=�l"�z	B9�ƪճ��S�02ŤHM�%���Q�wtiRE�a11�_�(����<�������C����e�,�	�1%�Y��)s�����?��%(���'��24�	1'L�d<o�#�U�u�WT�:&a:j��;�Jj�xa�ݽ9R�_X.;fV}P�"A���r��g����1��h�	1a�{cY����5����Z*5()�
շ��s�*-�F]���d�IW3���ժ��J��/u8�*i� w�q�/��܊�؋W���07"O�	�nA���=�s1<m
R���Pu�B���Pgu�7���vUY��%��b��6'�yx2AY���h~�x��˷�G ��q��$���#-V�;��e���Ăl�ˉo%ݒY ��s5�hA
j�lش=_���ާ��-)�CEUm�	Q�՘��{�R��3&����;z`r��'>3]R%l9X�[��3?��I�Q0��]B����
G�Q��[
G�i�?��Cؖ�k�,@
R�K����ʏ��$_�e���d��@ՙl�jS���n�Y��R�9�M�v8n��M��x���c^���P�Rˢжٛ �gzx����zg���K�W�9�:�o�ڔQϸ��3<)+yX�����p��qd��`��;q�E�9i3�� �l'A�ۀ��J�y�i|���/AmC�\UZ�܍Du�#0[��A����N5R{.��bh�s�D:ߪ�����'�*-	�:�ж�zH�+��E����C�P�U'pkː��E�x8w��m"uj6q�	��R��7&}r�c$��E�(G�]������j��u��)�o�NO
C�ňz�GKq�������0���ʎ)aɶ�.Q��S�'AU�E��LS�,�J�X�Ӓu��@�{�P=0N#WW�|�Zк`��X�+I\��4<�jL��j=\m���0LV'�/����w��    IEND�B`�PK
     �J�ZP��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     �J�Z$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK 
     �J�Z���sQ  sQ                   cirkitFile.jsonPK 
     �J�Z                        �Q  jsons/PK 
     �J�Z�haZ                 �Q  jsons/user_defined.jsonPK 
     �J�Z                        f  images/PK 
     �J�Z[�\� \� /             7f  images/707f98a2-ba92-4472-bb4e-3eede8d3998f.pngPK 
     �J�Z^R�#  �#  /             �3 images/e96e51a4-2e0a-4cc5-ba63-cf190e1d4d54.pngPK 
     �J�ZP��/ǽ  ǽ  /             �W images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     �J�Z$7h�!  �!  /             � images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK      _  %8   